module PositFMA31_3(
  input         clock,
  input         reset,
  input         io_inValid,
  input  [1:0]  io_fmaOp,
  input  [30:0] io_A,
  input  [30:0] io_B,
  input  [30:0] io_C,
  output [30:0] io_F,
  output        io_outValid
);
  wire  _T; // @[PositFMA.scala 47:36]
  wire [30:0] _T_2; // @[Bitwise.scala 71:12]
  wire [30:0] _T_3; // @[PositFMA.scala 47:41]
  wire [30:0] _GEN_10; // @[PositFMA.scala 47:49]
  wire [30:0] realA; // @[PositFMA.scala 47:49]
  wire  _T_6; // @[PositFMA.scala 48:36]
  wire [30:0] _T_8; // @[Bitwise.scala 71:12]
  wire [30:0] _T_9; // @[PositFMA.scala 48:41]
  wire [30:0] _GEN_11; // @[PositFMA.scala 48:49]
  wire [30:0] realC; // @[PositFMA.scala 48:49]
  wire  _T_13; // @[convert.scala 18:24]
  wire  _T_14; // @[convert.scala 18:40]
  wire  _T_15; // @[convert.scala 18:36]
  wire [28:0] _T_16; // @[convert.scala 19:24]
  wire [28:0] _T_17; // @[convert.scala 19:43]
  wire [28:0] _T_18; // @[convert.scala 19:39]
  wire [15:0] _T_19; // @[LZD.scala 43:32]
  wire [7:0] _T_20; // @[LZD.scala 43:32]
  wire [3:0] _T_21; // @[LZD.scala 43:32]
  wire [1:0] _T_22; // @[LZD.scala 43:32]
  wire  _T_23; // @[LZD.scala 39:14]
  wire  _T_24; // @[LZD.scala 39:21]
  wire  _T_25; // @[LZD.scala 39:30]
  wire  _T_26; // @[LZD.scala 39:27]
  wire  _T_27; // @[LZD.scala 39:25]
  wire [1:0] _T_28; // @[Cat.scala 29:58]
  wire [1:0] _T_29; // @[LZD.scala 44:32]
  wire  _T_30; // @[LZD.scala 39:14]
  wire  _T_31; // @[LZD.scala 39:21]
  wire  _T_32; // @[LZD.scala 39:30]
  wire  _T_33; // @[LZD.scala 39:27]
  wire  _T_34; // @[LZD.scala 39:25]
  wire [1:0] _T_35; // @[Cat.scala 29:58]
  wire  _T_36; // @[Shift.scala 12:21]
  wire  _T_37; // @[Shift.scala 12:21]
  wire  _T_38; // @[LZD.scala 49:16]
  wire  _T_39; // @[LZD.scala 49:27]
  wire  _T_40; // @[LZD.scala 49:25]
  wire  _T_41; // @[LZD.scala 49:47]
  wire  _T_42; // @[LZD.scala 49:59]
  wire  _T_43; // @[LZD.scala 49:35]
  wire [2:0] _T_45; // @[Cat.scala 29:58]
  wire [3:0] _T_46; // @[LZD.scala 44:32]
  wire [1:0] _T_47; // @[LZD.scala 43:32]
  wire  _T_48; // @[LZD.scala 39:14]
  wire  _T_49; // @[LZD.scala 39:21]
  wire  _T_50; // @[LZD.scala 39:30]
  wire  _T_51; // @[LZD.scala 39:27]
  wire  _T_52; // @[LZD.scala 39:25]
  wire [1:0] _T_53; // @[Cat.scala 29:58]
  wire [1:0] _T_54; // @[LZD.scala 44:32]
  wire  _T_55; // @[LZD.scala 39:14]
  wire  _T_56; // @[LZD.scala 39:21]
  wire  _T_57; // @[LZD.scala 39:30]
  wire  _T_58; // @[LZD.scala 39:27]
  wire  _T_59; // @[LZD.scala 39:25]
  wire [1:0] _T_60; // @[Cat.scala 29:58]
  wire  _T_61; // @[Shift.scala 12:21]
  wire  _T_62; // @[Shift.scala 12:21]
  wire  _T_63; // @[LZD.scala 49:16]
  wire  _T_64; // @[LZD.scala 49:27]
  wire  _T_65; // @[LZD.scala 49:25]
  wire  _T_66; // @[LZD.scala 49:47]
  wire  _T_67; // @[LZD.scala 49:59]
  wire  _T_68; // @[LZD.scala 49:35]
  wire [2:0] _T_70; // @[Cat.scala 29:58]
  wire  _T_71; // @[Shift.scala 12:21]
  wire  _T_72; // @[Shift.scala 12:21]
  wire  _T_73; // @[LZD.scala 49:16]
  wire  _T_74; // @[LZD.scala 49:27]
  wire  _T_75; // @[LZD.scala 49:25]
  wire [1:0] _T_76; // @[LZD.scala 49:47]
  wire [1:0] _T_77; // @[LZD.scala 49:59]
  wire [1:0] _T_78; // @[LZD.scala 49:35]
  wire [3:0] _T_80; // @[Cat.scala 29:58]
  wire [7:0] _T_81; // @[LZD.scala 44:32]
  wire [3:0] _T_82; // @[LZD.scala 43:32]
  wire [1:0] _T_83; // @[LZD.scala 43:32]
  wire  _T_84; // @[LZD.scala 39:14]
  wire  _T_85; // @[LZD.scala 39:21]
  wire  _T_86; // @[LZD.scala 39:30]
  wire  _T_87; // @[LZD.scala 39:27]
  wire  _T_88; // @[LZD.scala 39:25]
  wire [1:0] _T_89; // @[Cat.scala 29:58]
  wire [1:0] _T_90; // @[LZD.scala 44:32]
  wire  _T_91; // @[LZD.scala 39:14]
  wire  _T_92; // @[LZD.scala 39:21]
  wire  _T_93; // @[LZD.scala 39:30]
  wire  _T_94; // @[LZD.scala 39:27]
  wire  _T_95; // @[LZD.scala 39:25]
  wire [1:0] _T_96; // @[Cat.scala 29:58]
  wire  _T_97; // @[Shift.scala 12:21]
  wire  _T_98; // @[Shift.scala 12:21]
  wire  _T_99; // @[LZD.scala 49:16]
  wire  _T_100; // @[LZD.scala 49:27]
  wire  _T_101; // @[LZD.scala 49:25]
  wire  _T_102; // @[LZD.scala 49:47]
  wire  _T_103; // @[LZD.scala 49:59]
  wire  _T_104; // @[LZD.scala 49:35]
  wire [2:0] _T_106; // @[Cat.scala 29:58]
  wire [3:0] _T_107; // @[LZD.scala 44:32]
  wire [1:0] _T_108; // @[LZD.scala 43:32]
  wire  _T_109; // @[LZD.scala 39:14]
  wire  _T_110; // @[LZD.scala 39:21]
  wire  _T_111; // @[LZD.scala 39:30]
  wire  _T_112; // @[LZD.scala 39:27]
  wire  _T_113; // @[LZD.scala 39:25]
  wire [1:0] _T_114; // @[Cat.scala 29:58]
  wire [1:0] _T_115; // @[LZD.scala 44:32]
  wire  _T_116; // @[LZD.scala 39:14]
  wire  _T_117; // @[LZD.scala 39:21]
  wire  _T_118; // @[LZD.scala 39:30]
  wire  _T_119; // @[LZD.scala 39:27]
  wire  _T_120; // @[LZD.scala 39:25]
  wire [1:0] _T_121; // @[Cat.scala 29:58]
  wire  _T_122; // @[Shift.scala 12:21]
  wire  _T_123; // @[Shift.scala 12:21]
  wire  _T_124; // @[LZD.scala 49:16]
  wire  _T_125; // @[LZD.scala 49:27]
  wire  _T_126; // @[LZD.scala 49:25]
  wire  _T_127; // @[LZD.scala 49:47]
  wire  _T_128; // @[LZD.scala 49:59]
  wire  _T_129; // @[LZD.scala 49:35]
  wire [2:0] _T_131; // @[Cat.scala 29:58]
  wire  _T_132; // @[Shift.scala 12:21]
  wire  _T_133; // @[Shift.scala 12:21]
  wire  _T_134; // @[LZD.scala 49:16]
  wire  _T_135; // @[LZD.scala 49:27]
  wire  _T_136; // @[LZD.scala 49:25]
  wire [1:0] _T_137; // @[LZD.scala 49:47]
  wire [1:0] _T_138; // @[LZD.scala 49:59]
  wire [1:0] _T_139; // @[LZD.scala 49:35]
  wire [3:0] _T_141; // @[Cat.scala 29:58]
  wire  _T_142; // @[Shift.scala 12:21]
  wire  _T_143; // @[Shift.scala 12:21]
  wire  _T_144; // @[LZD.scala 49:16]
  wire  _T_145; // @[LZD.scala 49:27]
  wire  _T_146; // @[LZD.scala 49:25]
  wire [2:0] _T_147; // @[LZD.scala 49:47]
  wire [2:0] _T_148; // @[LZD.scala 49:59]
  wire [2:0] _T_149; // @[LZD.scala 49:35]
  wire [4:0] _T_151; // @[Cat.scala 29:58]
  wire [12:0] _T_152; // @[LZD.scala 44:32]
  wire [7:0] _T_153; // @[LZD.scala 43:32]
  wire [3:0] _T_154; // @[LZD.scala 43:32]
  wire [1:0] _T_155; // @[LZD.scala 43:32]
  wire  _T_156; // @[LZD.scala 39:14]
  wire  _T_157; // @[LZD.scala 39:21]
  wire  _T_158; // @[LZD.scala 39:30]
  wire  _T_159; // @[LZD.scala 39:27]
  wire  _T_160; // @[LZD.scala 39:25]
  wire [1:0] _T_161; // @[Cat.scala 29:58]
  wire [1:0] _T_162; // @[LZD.scala 44:32]
  wire  _T_163; // @[LZD.scala 39:14]
  wire  _T_164; // @[LZD.scala 39:21]
  wire  _T_165; // @[LZD.scala 39:30]
  wire  _T_166; // @[LZD.scala 39:27]
  wire  _T_167; // @[LZD.scala 39:25]
  wire [1:0] _T_168; // @[Cat.scala 29:58]
  wire  _T_169; // @[Shift.scala 12:21]
  wire  _T_170; // @[Shift.scala 12:21]
  wire  _T_171; // @[LZD.scala 49:16]
  wire  _T_172; // @[LZD.scala 49:27]
  wire  _T_173; // @[LZD.scala 49:25]
  wire  _T_174; // @[LZD.scala 49:47]
  wire  _T_175; // @[LZD.scala 49:59]
  wire  _T_176; // @[LZD.scala 49:35]
  wire [2:0] _T_178; // @[Cat.scala 29:58]
  wire [3:0] _T_179; // @[LZD.scala 44:32]
  wire [1:0] _T_180; // @[LZD.scala 43:32]
  wire  _T_181; // @[LZD.scala 39:14]
  wire  _T_182; // @[LZD.scala 39:21]
  wire  _T_183; // @[LZD.scala 39:30]
  wire  _T_184; // @[LZD.scala 39:27]
  wire  _T_185; // @[LZD.scala 39:25]
  wire [1:0] _T_186; // @[Cat.scala 29:58]
  wire [1:0] _T_187; // @[LZD.scala 44:32]
  wire  _T_188; // @[LZD.scala 39:14]
  wire  _T_189; // @[LZD.scala 39:21]
  wire  _T_190; // @[LZD.scala 39:30]
  wire  _T_191; // @[LZD.scala 39:27]
  wire  _T_192; // @[LZD.scala 39:25]
  wire [1:0] _T_193; // @[Cat.scala 29:58]
  wire  _T_194; // @[Shift.scala 12:21]
  wire  _T_195; // @[Shift.scala 12:21]
  wire  _T_196; // @[LZD.scala 49:16]
  wire  _T_197; // @[LZD.scala 49:27]
  wire  _T_198; // @[LZD.scala 49:25]
  wire  _T_199; // @[LZD.scala 49:47]
  wire  _T_200; // @[LZD.scala 49:59]
  wire  _T_201; // @[LZD.scala 49:35]
  wire [2:0] _T_203; // @[Cat.scala 29:58]
  wire  _T_204; // @[Shift.scala 12:21]
  wire  _T_205; // @[Shift.scala 12:21]
  wire  _T_206; // @[LZD.scala 49:16]
  wire  _T_207; // @[LZD.scala 49:27]
  wire  _T_208; // @[LZD.scala 49:25]
  wire [1:0] _T_209; // @[LZD.scala 49:47]
  wire [1:0] _T_210; // @[LZD.scala 49:59]
  wire [1:0] _T_211; // @[LZD.scala 49:35]
  wire [3:0] _T_213; // @[Cat.scala 29:58]
  wire [4:0] _T_214; // @[LZD.scala 44:32]
  wire [3:0] _T_215; // @[LZD.scala 43:32]
  wire [1:0] _T_216; // @[LZD.scala 43:32]
  wire  _T_217; // @[LZD.scala 39:14]
  wire  _T_218; // @[LZD.scala 39:21]
  wire  _T_219; // @[LZD.scala 39:30]
  wire  _T_220; // @[LZD.scala 39:27]
  wire  _T_221; // @[LZD.scala 39:25]
  wire [1:0] _T_222; // @[Cat.scala 29:58]
  wire [1:0] _T_223; // @[LZD.scala 44:32]
  wire  _T_224; // @[LZD.scala 39:14]
  wire  _T_225; // @[LZD.scala 39:21]
  wire  _T_226; // @[LZD.scala 39:30]
  wire  _T_227; // @[LZD.scala 39:27]
  wire  _T_228; // @[LZD.scala 39:25]
  wire [1:0] _T_229; // @[Cat.scala 29:58]
  wire  _T_230; // @[Shift.scala 12:21]
  wire  _T_231; // @[Shift.scala 12:21]
  wire  _T_232; // @[LZD.scala 49:16]
  wire  _T_233; // @[LZD.scala 49:27]
  wire  _T_234; // @[LZD.scala 49:25]
  wire  _T_235; // @[LZD.scala 49:47]
  wire  _T_236; // @[LZD.scala 49:59]
  wire  _T_237; // @[LZD.scala 49:35]
  wire [2:0] _T_239; // @[Cat.scala 29:58]
  wire  _T_240; // @[LZD.scala 44:32]
  wire  _T_242; // @[Shift.scala 12:21]
  wire [1:0] _T_244; // @[Cat.scala 29:58]
  wire [1:0] _T_245; // @[LZD.scala 55:32]
  wire [1:0] _T_246; // @[LZD.scala 55:20]
  wire [2:0] _T_247; // @[Cat.scala 29:58]
  wire  _T_248; // @[Shift.scala 12:21]
  wire [2:0] _T_250; // @[LZD.scala 55:32]
  wire [2:0] _T_251; // @[LZD.scala 55:20]
  wire [3:0] _T_252; // @[Cat.scala 29:58]
  wire  _T_253; // @[Shift.scala 12:21]
  wire [3:0] _T_255; // @[LZD.scala 55:32]
  wire [3:0] _T_256; // @[LZD.scala 55:20]
  wire [4:0] _T_257; // @[Cat.scala 29:58]
  wire [4:0] _T_258; // @[convert.scala 21:22]
  wire [27:0] _T_259; // @[convert.scala 22:36]
  wire  _T_260; // @[Shift.scala 16:24]
  wire  _T_262; // @[Shift.scala 12:21]
  wire [11:0] _T_263; // @[Shift.scala 64:52]
  wire [27:0] _T_265; // @[Cat.scala 29:58]
  wire [27:0] _T_266; // @[Shift.scala 64:27]
  wire [3:0] _T_267; // @[Shift.scala 66:70]
  wire  _T_268; // @[Shift.scala 12:21]
  wire [19:0] _T_269; // @[Shift.scala 64:52]
  wire [27:0] _T_271; // @[Cat.scala 29:58]
  wire [27:0] _T_272; // @[Shift.scala 64:27]
  wire [2:0] _T_273; // @[Shift.scala 66:70]
  wire  _T_274; // @[Shift.scala 12:21]
  wire [23:0] _T_275; // @[Shift.scala 64:52]
  wire [27:0] _T_277; // @[Cat.scala 29:58]
  wire [27:0] _T_278; // @[Shift.scala 64:27]
  wire [1:0] _T_279; // @[Shift.scala 66:70]
  wire  _T_280; // @[Shift.scala 12:21]
  wire [25:0] _T_281; // @[Shift.scala 64:52]
  wire [27:0] _T_283; // @[Cat.scala 29:58]
  wire [27:0] _T_284; // @[Shift.scala 64:27]
  wire  _T_285; // @[Shift.scala 66:70]
  wire [26:0] _T_287; // @[Shift.scala 64:52]
  wire [27:0] _T_288; // @[Cat.scala 29:58]
  wire [27:0] _T_289; // @[Shift.scala 64:27]
  wire [27:0] _T_290; // @[Shift.scala 16:10]
  wire [2:0] _T_291; // @[convert.scala 23:34]
  wire [24:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_293; // @[convert.scala 25:26]
  wire [4:0] _T_295; // @[convert.scala 25:42]
  wire [2:0] _T_298; // @[convert.scala 26:67]
  wire [2:0] _T_299; // @[convert.scala 26:51]
  wire [8:0] _T_300; // @[Cat.scala 29:58]
  wire [29:0] _T_302; // @[convert.scala 29:56]
  wire  _T_303; // @[convert.scala 29:60]
  wire  _T_304; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_307; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [8:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_316; // @[convert.scala 18:24]
  wire  _T_317; // @[convert.scala 18:40]
  wire  _T_318; // @[convert.scala 18:36]
  wire [28:0] _T_319; // @[convert.scala 19:24]
  wire [28:0] _T_320; // @[convert.scala 19:43]
  wire [28:0] _T_321; // @[convert.scala 19:39]
  wire [15:0] _T_322; // @[LZD.scala 43:32]
  wire [7:0] _T_323; // @[LZD.scala 43:32]
  wire [3:0] _T_324; // @[LZD.scala 43:32]
  wire [1:0] _T_325; // @[LZD.scala 43:32]
  wire  _T_326; // @[LZD.scala 39:14]
  wire  _T_327; // @[LZD.scala 39:21]
  wire  _T_328; // @[LZD.scala 39:30]
  wire  _T_329; // @[LZD.scala 39:27]
  wire  _T_330; // @[LZD.scala 39:25]
  wire [1:0] _T_331; // @[Cat.scala 29:58]
  wire [1:0] _T_332; // @[LZD.scala 44:32]
  wire  _T_333; // @[LZD.scala 39:14]
  wire  _T_334; // @[LZD.scala 39:21]
  wire  _T_335; // @[LZD.scala 39:30]
  wire  _T_336; // @[LZD.scala 39:27]
  wire  _T_337; // @[LZD.scala 39:25]
  wire [1:0] _T_338; // @[Cat.scala 29:58]
  wire  _T_339; // @[Shift.scala 12:21]
  wire  _T_340; // @[Shift.scala 12:21]
  wire  _T_341; // @[LZD.scala 49:16]
  wire  _T_342; // @[LZD.scala 49:27]
  wire  _T_343; // @[LZD.scala 49:25]
  wire  _T_344; // @[LZD.scala 49:47]
  wire  _T_345; // @[LZD.scala 49:59]
  wire  _T_346; // @[LZD.scala 49:35]
  wire [2:0] _T_348; // @[Cat.scala 29:58]
  wire [3:0] _T_349; // @[LZD.scala 44:32]
  wire [1:0] _T_350; // @[LZD.scala 43:32]
  wire  _T_351; // @[LZD.scala 39:14]
  wire  _T_352; // @[LZD.scala 39:21]
  wire  _T_353; // @[LZD.scala 39:30]
  wire  _T_354; // @[LZD.scala 39:27]
  wire  _T_355; // @[LZD.scala 39:25]
  wire [1:0] _T_356; // @[Cat.scala 29:58]
  wire [1:0] _T_357; // @[LZD.scala 44:32]
  wire  _T_358; // @[LZD.scala 39:14]
  wire  _T_359; // @[LZD.scala 39:21]
  wire  _T_360; // @[LZD.scala 39:30]
  wire  _T_361; // @[LZD.scala 39:27]
  wire  _T_362; // @[LZD.scala 39:25]
  wire [1:0] _T_363; // @[Cat.scala 29:58]
  wire  _T_364; // @[Shift.scala 12:21]
  wire  _T_365; // @[Shift.scala 12:21]
  wire  _T_366; // @[LZD.scala 49:16]
  wire  _T_367; // @[LZD.scala 49:27]
  wire  _T_368; // @[LZD.scala 49:25]
  wire  _T_369; // @[LZD.scala 49:47]
  wire  _T_370; // @[LZD.scala 49:59]
  wire  _T_371; // @[LZD.scala 49:35]
  wire [2:0] _T_373; // @[Cat.scala 29:58]
  wire  _T_374; // @[Shift.scala 12:21]
  wire  _T_375; // @[Shift.scala 12:21]
  wire  _T_376; // @[LZD.scala 49:16]
  wire  _T_377; // @[LZD.scala 49:27]
  wire  _T_378; // @[LZD.scala 49:25]
  wire [1:0] _T_379; // @[LZD.scala 49:47]
  wire [1:0] _T_380; // @[LZD.scala 49:59]
  wire [1:0] _T_381; // @[LZD.scala 49:35]
  wire [3:0] _T_383; // @[Cat.scala 29:58]
  wire [7:0] _T_384; // @[LZD.scala 44:32]
  wire [3:0] _T_385; // @[LZD.scala 43:32]
  wire [1:0] _T_386; // @[LZD.scala 43:32]
  wire  _T_387; // @[LZD.scala 39:14]
  wire  _T_388; // @[LZD.scala 39:21]
  wire  _T_389; // @[LZD.scala 39:30]
  wire  _T_390; // @[LZD.scala 39:27]
  wire  _T_391; // @[LZD.scala 39:25]
  wire [1:0] _T_392; // @[Cat.scala 29:58]
  wire [1:0] _T_393; // @[LZD.scala 44:32]
  wire  _T_394; // @[LZD.scala 39:14]
  wire  _T_395; // @[LZD.scala 39:21]
  wire  _T_396; // @[LZD.scala 39:30]
  wire  _T_397; // @[LZD.scala 39:27]
  wire  _T_398; // @[LZD.scala 39:25]
  wire [1:0] _T_399; // @[Cat.scala 29:58]
  wire  _T_400; // @[Shift.scala 12:21]
  wire  _T_401; // @[Shift.scala 12:21]
  wire  _T_402; // @[LZD.scala 49:16]
  wire  _T_403; // @[LZD.scala 49:27]
  wire  _T_404; // @[LZD.scala 49:25]
  wire  _T_405; // @[LZD.scala 49:47]
  wire  _T_406; // @[LZD.scala 49:59]
  wire  _T_407; // @[LZD.scala 49:35]
  wire [2:0] _T_409; // @[Cat.scala 29:58]
  wire [3:0] _T_410; // @[LZD.scala 44:32]
  wire [1:0] _T_411; // @[LZD.scala 43:32]
  wire  _T_412; // @[LZD.scala 39:14]
  wire  _T_413; // @[LZD.scala 39:21]
  wire  _T_414; // @[LZD.scala 39:30]
  wire  _T_415; // @[LZD.scala 39:27]
  wire  _T_416; // @[LZD.scala 39:25]
  wire [1:0] _T_417; // @[Cat.scala 29:58]
  wire [1:0] _T_418; // @[LZD.scala 44:32]
  wire  _T_419; // @[LZD.scala 39:14]
  wire  _T_420; // @[LZD.scala 39:21]
  wire  _T_421; // @[LZD.scala 39:30]
  wire  _T_422; // @[LZD.scala 39:27]
  wire  _T_423; // @[LZD.scala 39:25]
  wire [1:0] _T_424; // @[Cat.scala 29:58]
  wire  _T_425; // @[Shift.scala 12:21]
  wire  _T_426; // @[Shift.scala 12:21]
  wire  _T_427; // @[LZD.scala 49:16]
  wire  _T_428; // @[LZD.scala 49:27]
  wire  _T_429; // @[LZD.scala 49:25]
  wire  _T_430; // @[LZD.scala 49:47]
  wire  _T_431; // @[LZD.scala 49:59]
  wire  _T_432; // @[LZD.scala 49:35]
  wire [2:0] _T_434; // @[Cat.scala 29:58]
  wire  _T_435; // @[Shift.scala 12:21]
  wire  _T_436; // @[Shift.scala 12:21]
  wire  _T_437; // @[LZD.scala 49:16]
  wire  _T_438; // @[LZD.scala 49:27]
  wire  _T_439; // @[LZD.scala 49:25]
  wire [1:0] _T_440; // @[LZD.scala 49:47]
  wire [1:0] _T_441; // @[LZD.scala 49:59]
  wire [1:0] _T_442; // @[LZD.scala 49:35]
  wire [3:0] _T_444; // @[Cat.scala 29:58]
  wire  _T_445; // @[Shift.scala 12:21]
  wire  _T_446; // @[Shift.scala 12:21]
  wire  _T_447; // @[LZD.scala 49:16]
  wire  _T_448; // @[LZD.scala 49:27]
  wire  _T_449; // @[LZD.scala 49:25]
  wire [2:0] _T_450; // @[LZD.scala 49:47]
  wire [2:0] _T_451; // @[LZD.scala 49:59]
  wire [2:0] _T_452; // @[LZD.scala 49:35]
  wire [4:0] _T_454; // @[Cat.scala 29:58]
  wire [12:0] _T_455; // @[LZD.scala 44:32]
  wire [7:0] _T_456; // @[LZD.scala 43:32]
  wire [3:0] _T_457; // @[LZD.scala 43:32]
  wire [1:0] _T_458; // @[LZD.scala 43:32]
  wire  _T_459; // @[LZD.scala 39:14]
  wire  _T_460; // @[LZD.scala 39:21]
  wire  _T_461; // @[LZD.scala 39:30]
  wire  _T_462; // @[LZD.scala 39:27]
  wire  _T_463; // @[LZD.scala 39:25]
  wire [1:0] _T_464; // @[Cat.scala 29:58]
  wire [1:0] _T_465; // @[LZD.scala 44:32]
  wire  _T_466; // @[LZD.scala 39:14]
  wire  _T_467; // @[LZD.scala 39:21]
  wire  _T_468; // @[LZD.scala 39:30]
  wire  _T_469; // @[LZD.scala 39:27]
  wire  _T_470; // @[LZD.scala 39:25]
  wire [1:0] _T_471; // @[Cat.scala 29:58]
  wire  _T_472; // @[Shift.scala 12:21]
  wire  _T_473; // @[Shift.scala 12:21]
  wire  _T_474; // @[LZD.scala 49:16]
  wire  _T_475; // @[LZD.scala 49:27]
  wire  _T_476; // @[LZD.scala 49:25]
  wire  _T_477; // @[LZD.scala 49:47]
  wire  _T_478; // @[LZD.scala 49:59]
  wire  _T_479; // @[LZD.scala 49:35]
  wire [2:0] _T_481; // @[Cat.scala 29:58]
  wire [3:0] _T_482; // @[LZD.scala 44:32]
  wire [1:0] _T_483; // @[LZD.scala 43:32]
  wire  _T_484; // @[LZD.scala 39:14]
  wire  _T_485; // @[LZD.scala 39:21]
  wire  _T_486; // @[LZD.scala 39:30]
  wire  _T_487; // @[LZD.scala 39:27]
  wire  _T_488; // @[LZD.scala 39:25]
  wire [1:0] _T_489; // @[Cat.scala 29:58]
  wire [1:0] _T_490; // @[LZD.scala 44:32]
  wire  _T_491; // @[LZD.scala 39:14]
  wire  _T_492; // @[LZD.scala 39:21]
  wire  _T_493; // @[LZD.scala 39:30]
  wire  _T_494; // @[LZD.scala 39:27]
  wire  _T_495; // @[LZD.scala 39:25]
  wire [1:0] _T_496; // @[Cat.scala 29:58]
  wire  _T_497; // @[Shift.scala 12:21]
  wire  _T_498; // @[Shift.scala 12:21]
  wire  _T_499; // @[LZD.scala 49:16]
  wire  _T_500; // @[LZD.scala 49:27]
  wire  _T_501; // @[LZD.scala 49:25]
  wire  _T_502; // @[LZD.scala 49:47]
  wire  _T_503; // @[LZD.scala 49:59]
  wire  _T_504; // @[LZD.scala 49:35]
  wire [2:0] _T_506; // @[Cat.scala 29:58]
  wire  _T_507; // @[Shift.scala 12:21]
  wire  _T_508; // @[Shift.scala 12:21]
  wire  _T_509; // @[LZD.scala 49:16]
  wire  _T_510; // @[LZD.scala 49:27]
  wire  _T_511; // @[LZD.scala 49:25]
  wire [1:0] _T_512; // @[LZD.scala 49:47]
  wire [1:0] _T_513; // @[LZD.scala 49:59]
  wire [1:0] _T_514; // @[LZD.scala 49:35]
  wire [3:0] _T_516; // @[Cat.scala 29:58]
  wire [4:0] _T_517; // @[LZD.scala 44:32]
  wire [3:0] _T_518; // @[LZD.scala 43:32]
  wire [1:0] _T_519; // @[LZD.scala 43:32]
  wire  _T_520; // @[LZD.scala 39:14]
  wire  _T_521; // @[LZD.scala 39:21]
  wire  _T_522; // @[LZD.scala 39:30]
  wire  _T_523; // @[LZD.scala 39:27]
  wire  _T_524; // @[LZD.scala 39:25]
  wire [1:0] _T_525; // @[Cat.scala 29:58]
  wire [1:0] _T_526; // @[LZD.scala 44:32]
  wire  _T_527; // @[LZD.scala 39:14]
  wire  _T_528; // @[LZD.scala 39:21]
  wire  _T_529; // @[LZD.scala 39:30]
  wire  _T_530; // @[LZD.scala 39:27]
  wire  _T_531; // @[LZD.scala 39:25]
  wire [1:0] _T_532; // @[Cat.scala 29:58]
  wire  _T_533; // @[Shift.scala 12:21]
  wire  _T_534; // @[Shift.scala 12:21]
  wire  _T_535; // @[LZD.scala 49:16]
  wire  _T_536; // @[LZD.scala 49:27]
  wire  _T_537; // @[LZD.scala 49:25]
  wire  _T_538; // @[LZD.scala 49:47]
  wire  _T_539; // @[LZD.scala 49:59]
  wire  _T_540; // @[LZD.scala 49:35]
  wire [2:0] _T_542; // @[Cat.scala 29:58]
  wire  _T_543; // @[LZD.scala 44:32]
  wire  _T_545; // @[Shift.scala 12:21]
  wire [1:0] _T_547; // @[Cat.scala 29:58]
  wire [1:0] _T_548; // @[LZD.scala 55:32]
  wire [1:0] _T_549; // @[LZD.scala 55:20]
  wire [2:0] _T_550; // @[Cat.scala 29:58]
  wire  _T_551; // @[Shift.scala 12:21]
  wire [2:0] _T_553; // @[LZD.scala 55:32]
  wire [2:0] _T_554; // @[LZD.scala 55:20]
  wire [3:0] _T_555; // @[Cat.scala 29:58]
  wire  _T_556; // @[Shift.scala 12:21]
  wire [3:0] _T_558; // @[LZD.scala 55:32]
  wire [3:0] _T_559; // @[LZD.scala 55:20]
  wire [4:0] _T_560; // @[Cat.scala 29:58]
  wire [4:0] _T_561; // @[convert.scala 21:22]
  wire [27:0] _T_562; // @[convert.scala 22:36]
  wire  _T_563; // @[Shift.scala 16:24]
  wire  _T_565; // @[Shift.scala 12:21]
  wire [11:0] _T_566; // @[Shift.scala 64:52]
  wire [27:0] _T_568; // @[Cat.scala 29:58]
  wire [27:0] _T_569; // @[Shift.scala 64:27]
  wire [3:0] _T_570; // @[Shift.scala 66:70]
  wire  _T_571; // @[Shift.scala 12:21]
  wire [19:0] _T_572; // @[Shift.scala 64:52]
  wire [27:0] _T_574; // @[Cat.scala 29:58]
  wire [27:0] _T_575; // @[Shift.scala 64:27]
  wire [2:0] _T_576; // @[Shift.scala 66:70]
  wire  _T_577; // @[Shift.scala 12:21]
  wire [23:0] _T_578; // @[Shift.scala 64:52]
  wire [27:0] _T_580; // @[Cat.scala 29:58]
  wire [27:0] _T_581; // @[Shift.scala 64:27]
  wire [1:0] _T_582; // @[Shift.scala 66:70]
  wire  _T_583; // @[Shift.scala 12:21]
  wire [25:0] _T_584; // @[Shift.scala 64:52]
  wire [27:0] _T_586; // @[Cat.scala 29:58]
  wire [27:0] _T_587; // @[Shift.scala 64:27]
  wire  _T_588; // @[Shift.scala 66:70]
  wire [26:0] _T_590; // @[Shift.scala 64:52]
  wire [27:0] _T_591; // @[Cat.scala 29:58]
  wire [27:0] _T_592; // @[Shift.scala 64:27]
  wire [27:0] _T_593; // @[Shift.scala 16:10]
  wire [2:0] _T_594; // @[convert.scala 23:34]
  wire [24:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_596; // @[convert.scala 25:26]
  wire [4:0] _T_598; // @[convert.scala 25:42]
  wire [2:0] _T_601; // @[convert.scala 26:67]
  wire [2:0] _T_602; // @[convert.scala 26:51]
  wire [8:0] _T_603; // @[Cat.scala 29:58]
  wire [29:0] _T_605; // @[convert.scala 29:56]
  wire  _T_606; // @[convert.scala 29:60]
  wire  _T_607; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_610; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [8:0] decB_scale; // @[convert.scala 32:24]
  wire  _T_619; // @[convert.scala 18:24]
  wire  _T_620; // @[convert.scala 18:40]
  wire  _T_621; // @[convert.scala 18:36]
  wire [28:0] _T_622; // @[convert.scala 19:24]
  wire [28:0] _T_623; // @[convert.scala 19:43]
  wire [28:0] _T_624; // @[convert.scala 19:39]
  wire [15:0] _T_625; // @[LZD.scala 43:32]
  wire [7:0] _T_626; // @[LZD.scala 43:32]
  wire [3:0] _T_627; // @[LZD.scala 43:32]
  wire [1:0] _T_628; // @[LZD.scala 43:32]
  wire  _T_629; // @[LZD.scala 39:14]
  wire  _T_630; // @[LZD.scala 39:21]
  wire  _T_631; // @[LZD.scala 39:30]
  wire  _T_632; // @[LZD.scala 39:27]
  wire  _T_633; // @[LZD.scala 39:25]
  wire [1:0] _T_634; // @[Cat.scala 29:58]
  wire [1:0] _T_635; // @[LZD.scala 44:32]
  wire  _T_636; // @[LZD.scala 39:14]
  wire  _T_637; // @[LZD.scala 39:21]
  wire  _T_638; // @[LZD.scala 39:30]
  wire  _T_639; // @[LZD.scala 39:27]
  wire  _T_640; // @[LZD.scala 39:25]
  wire [1:0] _T_641; // @[Cat.scala 29:58]
  wire  _T_642; // @[Shift.scala 12:21]
  wire  _T_643; // @[Shift.scala 12:21]
  wire  _T_644; // @[LZD.scala 49:16]
  wire  _T_645; // @[LZD.scala 49:27]
  wire  _T_646; // @[LZD.scala 49:25]
  wire  _T_647; // @[LZD.scala 49:47]
  wire  _T_648; // @[LZD.scala 49:59]
  wire  _T_649; // @[LZD.scala 49:35]
  wire [2:0] _T_651; // @[Cat.scala 29:58]
  wire [3:0] _T_652; // @[LZD.scala 44:32]
  wire [1:0] _T_653; // @[LZD.scala 43:32]
  wire  _T_654; // @[LZD.scala 39:14]
  wire  _T_655; // @[LZD.scala 39:21]
  wire  _T_656; // @[LZD.scala 39:30]
  wire  _T_657; // @[LZD.scala 39:27]
  wire  _T_658; // @[LZD.scala 39:25]
  wire [1:0] _T_659; // @[Cat.scala 29:58]
  wire [1:0] _T_660; // @[LZD.scala 44:32]
  wire  _T_661; // @[LZD.scala 39:14]
  wire  _T_662; // @[LZD.scala 39:21]
  wire  _T_663; // @[LZD.scala 39:30]
  wire  _T_664; // @[LZD.scala 39:27]
  wire  _T_665; // @[LZD.scala 39:25]
  wire [1:0] _T_666; // @[Cat.scala 29:58]
  wire  _T_667; // @[Shift.scala 12:21]
  wire  _T_668; // @[Shift.scala 12:21]
  wire  _T_669; // @[LZD.scala 49:16]
  wire  _T_670; // @[LZD.scala 49:27]
  wire  _T_671; // @[LZD.scala 49:25]
  wire  _T_672; // @[LZD.scala 49:47]
  wire  _T_673; // @[LZD.scala 49:59]
  wire  _T_674; // @[LZD.scala 49:35]
  wire [2:0] _T_676; // @[Cat.scala 29:58]
  wire  _T_677; // @[Shift.scala 12:21]
  wire  _T_678; // @[Shift.scala 12:21]
  wire  _T_679; // @[LZD.scala 49:16]
  wire  _T_680; // @[LZD.scala 49:27]
  wire  _T_681; // @[LZD.scala 49:25]
  wire [1:0] _T_682; // @[LZD.scala 49:47]
  wire [1:0] _T_683; // @[LZD.scala 49:59]
  wire [1:0] _T_684; // @[LZD.scala 49:35]
  wire [3:0] _T_686; // @[Cat.scala 29:58]
  wire [7:0] _T_687; // @[LZD.scala 44:32]
  wire [3:0] _T_688; // @[LZD.scala 43:32]
  wire [1:0] _T_689; // @[LZD.scala 43:32]
  wire  _T_690; // @[LZD.scala 39:14]
  wire  _T_691; // @[LZD.scala 39:21]
  wire  _T_692; // @[LZD.scala 39:30]
  wire  _T_693; // @[LZD.scala 39:27]
  wire  _T_694; // @[LZD.scala 39:25]
  wire [1:0] _T_695; // @[Cat.scala 29:58]
  wire [1:0] _T_696; // @[LZD.scala 44:32]
  wire  _T_697; // @[LZD.scala 39:14]
  wire  _T_698; // @[LZD.scala 39:21]
  wire  _T_699; // @[LZD.scala 39:30]
  wire  _T_700; // @[LZD.scala 39:27]
  wire  _T_701; // @[LZD.scala 39:25]
  wire [1:0] _T_702; // @[Cat.scala 29:58]
  wire  _T_703; // @[Shift.scala 12:21]
  wire  _T_704; // @[Shift.scala 12:21]
  wire  _T_705; // @[LZD.scala 49:16]
  wire  _T_706; // @[LZD.scala 49:27]
  wire  _T_707; // @[LZD.scala 49:25]
  wire  _T_708; // @[LZD.scala 49:47]
  wire  _T_709; // @[LZD.scala 49:59]
  wire  _T_710; // @[LZD.scala 49:35]
  wire [2:0] _T_712; // @[Cat.scala 29:58]
  wire [3:0] _T_713; // @[LZD.scala 44:32]
  wire [1:0] _T_714; // @[LZD.scala 43:32]
  wire  _T_715; // @[LZD.scala 39:14]
  wire  _T_716; // @[LZD.scala 39:21]
  wire  _T_717; // @[LZD.scala 39:30]
  wire  _T_718; // @[LZD.scala 39:27]
  wire  _T_719; // @[LZD.scala 39:25]
  wire [1:0] _T_720; // @[Cat.scala 29:58]
  wire [1:0] _T_721; // @[LZD.scala 44:32]
  wire  _T_722; // @[LZD.scala 39:14]
  wire  _T_723; // @[LZD.scala 39:21]
  wire  _T_724; // @[LZD.scala 39:30]
  wire  _T_725; // @[LZD.scala 39:27]
  wire  _T_726; // @[LZD.scala 39:25]
  wire [1:0] _T_727; // @[Cat.scala 29:58]
  wire  _T_728; // @[Shift.scala 12:21]
  wire  _T_729; // @[Shift.scala 12:21]
  wire  _T_730; // @[LZD.scala 49:16]
  wire  _T_731; // @[LZD.scala 49:27]
  wire  _T_732; // @[LZD.scala 49:25]
  wire  _T_733; // @[LZD.scala 49:47]
  wire  _T_734; // @[LZD.scala 49:59]
  wire  _T_735; // @[LZD.scala 49:35]
  wire [2:0] _T_737; // @[Cat.scala 29:58]
  wire  _T_738; // @[Shift.scala 12:21]
  wire  _T_739; // @[Shift.scala 12:21]
  wire  _T_740; // @[LZD.scala 49:16]
  wire  _T_741; // @[LZD.scala 49:27]
  wire  _T_742; // @[LZD.scala 49:25]
  wire [1:0] _T_743; // @[LZD.scala 49:47]
  wire [1:0] _T_744; // @[LZD.scala 49:59]
  wire [1:0] _T_745; // @[LZD.scala 49:35]
  wire [3:0] _T_747; // @[Cat.scala 29:58]
  wire  _T_748; // @[Shift.scala 12:21]
  wire  _T_749; // @[Shift.scala 12:21]
  wire  _T_750; // @[LZD.scala 49:16]
  wire  _T_751; // @[LZD.scala 49:27]
  wire  _T_752; // @[LZD.scala 49:25]
  wire [2:0] _T_753; // @[LZD.scala 49:47]
  wire [2:0] _T_754; // @[LZD.scala 49:59]
  wire [2:0] _T_755; // @[LZD.scala 49:35]
  wire [4:0] _T_757; // @[Cat.scala 29:58]
  wire [12:0] _T_758; // @[LZD.scala 44:32]
  wire [7:0] _T_759; // @[LZD.scala 43:32]
  wire [3:0] _T_760; // @[LZD.scala 43:32]
  wire [1:0] _T_761; // @[LZD.scala 43:32]
  wire  _T_762; // @[LZD.scala 39:14]
  wire  _T_763; // @[LZD.scala 39:21]
  wire  _T_764; // @[LZD.scala 39:30]
  wire  _T_765; // @[LZD.scala 39:27]
  wire  _T_766; // @[LZD.scala 39:25]
  wire [1:0] _T_767; // @[Cat.scala 29:58]
  wire [1:0] _T_768; // @[LZD.scala 44:32]
  wire  _T_769; // @[LZD.scala 39:14]
  wire  _T_770; // @[LZD.scala 39:21]
  wire  _T_771; // @[LZD.scala 39:30]
  wire  _T_772; // @[LZD.scala 39:27]
  wire  _T_773; // @[LZD.scala 39:25]
  wire [1:0] _T_774; // @[Cat.scala 29:58]
  wire  _T_775; // @[Shift.scala 12:21]
  wire  _T_776; // @[Shift.scala 12:21]
  wire  _T_777; // @[LZD.scala 49:16]
  wire  _T_778; // @[LZD.scala 49:27]
  wire  _T_779; // @[LZD.scala 49:25]
  wire  _T_780; // @[LZD.scala 49:47]
  wire  _T_781; // @[LZD.scala 49:59]
  wire  _T_782; // @[LZD.scala 49:35]
  wire [2:0] _T_784; // @[Cat.scala 29:58]
  wire [3:0] _T_785; // @[LZD.scala 44:32]
  wire [1:0] _T_786; // @[LZD.scala 43:32]
  wire  _T_787; // @[LZD.scala 39:14]
  wire  _T_788; // @[LZD.scala 39:21]
  wire  _T_789; // @[LZD.scala 39:30]
  wire  _T_790; // @[LZD.scala 39:27]
  wire  _T_791; // @[LZD.scala 39:25]
  wire [1:0] _T_792; // @[Cat.scala 29:58]
  wire [1:0] _T_793; // @[LZD.scala 44:32]
  wire  _T_794; // @[LZD.scala 39:14]
  wire  _T_795; // @[LZD.scala 39:21]
  wire  _T_796; // @[LZD.scala 39:30]
  wire  _T_797; // @[LZD.scala 39:27]
  wire  _T_798; // @[LZD.scala 39:25]
  wire [1:0] _T_799; // @[Cat.scala 29:58]
  wire  _T_800; // @[Shift.scala 12:21]
  wire  _T_801; // @[Shift.scala 12:21]
  wire  _T_802; // @[LZD.scala 49:16]
  wire  _T_803; // @[LZD.scala 49:27]
  wire  _T_804; // @[LZD.scala 49:25]
  wire  _T_805; // @[LZD.scala 49:47]
  wire  _T_806; // @[LZD.scala 49:59]
  wire  _T_807; // @[LZD.scala 49:35]
  wire [2:0] _T_809; // @[Cat.scala 29:58]
  wire  _T_810; // @[Shift.scala 12:21]
  wire  _T_811; // @[Shift.scala 12:21]
  wire  _T_812; // @[LZD.scala 49:16]
  wire  _T_813; // @[LZD.scala 49:27]
  wire  _T_814; // @[LZD.scala 49:25]
  wire [1:0] _T_815; // @[LZD.scala 49:47]
  wire [1:0] _T_816; // @[LZD.scala 49:59]
  wire [1:0] _T_817; // @[LZD.scala 49:35]
  wire [3:0] _T_819; // @[Cat.scala 29:58]
  wire [4:0] _T_820; // @[LZD.scala 44:32]
  wire [3:0] _T_821; // @[LZD.scala 43:32]
  wire [1:0] _T_822; // @[LZD.scala 43:32]
  wire  _T_823; // @[LZD.scala 39:14]
  wire  _T_824; // @[LZD.scala 39:21]
  wire  _T_825; // @[LZD.scala 39:30]
  wire  _T_826; // @[LZD.scala 39:27]
  wire  _T_827; // @[LZD.scala 39:25]
  wire [1:0] _T_828; // @[Cat.scala 29:58]
  wire [1:0] _T_829; // @[LZD.scala 44:32]
  wire  _T_830; // @[LZD.scala 39:14]
  wire  _T_831; // @[LZD.scala 39:21]
  wire  _T_832; // @[LZD.scala 39:30]
  wire  _T_833; // @[LZD.scala 39:27]
  wire  _T_834; // @[LZD.scala 39:25]
  wire [1:0] _T_835; // @[Cat.scala 29:58]
  wire  _T_836; // @[Shift.scala 12:21]
  wire  _T_837; // @[Shift.scala 12:21]
  wire  _T_838; // @[LZD.scala 49:16]
  wire  _T_839; // @[LZD.scala 49:27]
  wire  _T_840; // @[LZD.scala 49:25]
  wire  _T_841; // @[LZD.scala 49:47]
  wire  _T_842; // @[LZD.scala 49:59]
  wire  _T_843; // @[LZD.scala 49:35]
  wire [2:0] _T_845; // @[Cat.scala 29:58]
  wire  _T_846; // @[LZD.scala 44:32]
  wire  _T_848; // @[Shift.scala 12:21]
  wire [1:0] _T_850; // @[Cat.scala 29:58]
  wire [1:0] _T_851; // @[LZD.scala 55:32]
  wire [1:0] _T_852; // @[LZD.scala 55:20]
  wire [2:0] _T_853; // @[Cat.scala 29:58]
  wire  _T_854; // @[Shift.scala 12:21]
  wire [2:0] _T_856; // @[LZD.scala 55:32]
  wire [2:0] _T_857; // @[LZD.scala 55:20]
  wire [3:0] _T_858; // @[Cat.scala 29:58]
  wire  _T_859; // @[Shift.scala 12:21]
  wire [3:0] _T_861; // @[LZD.scala 55:32]
  wire [3:0] _T_862; // @[LZD.scala 55:20]
  wire [4:0] _T_863; // @[Cat.scala 29:58]
  wire [4:0] _T_864; // @[convert.scala 21:22]
  wire [27:0] _T_865; // @[convert.scala 22:36]
  wire  _T_866; // @[Shift.scala 16:24]
  wire  _T_868; // @[Shift.scala 12:21]
  wire [11:0] _T_869; // @[Shift.scala 64:52]
  wire [27:0] _T_871; // @[Cat.scala 29:58]
  wire [27:0] _T_872; // @[Shift.scala 64:27]
  wire [3:0] _T_873; // @[Shift.scala 66:70]
  wire  _T_874; // @[Shift.scala 12:21]
  wire [19:0] _T_875; // @[Shift.scala 64:52]
  wire [27:0] _T_877; // @[Cat.scala 29:58]
  wire [27:0] _T_878; // @[Shift.scala 64:27]
  wire [2:0] _T_879; // @[Shift.scala 66:70]
  wire  _T_880; // @[Shift.scala 12:21]
  wire [23:0] _T_881; // @[Shift.scala 64:52]
  wire [27:0] _T_883; // @[Cat.scala 29:58]
  wire [27:0] _T_884; // @[Shift.scala 64:27]
  wire [1:0] _T_885; // @[Shift.scala 66:70]
  wire  _T_886; // @[Shift.scala 12:21]
  wire [25:0] _T_887; // @[Shift.scala 64:52]
  wire [27:0] _T_889; // @[Cat.scala 29:58]
  wire [27:0] _T_890; // @[Shift.scala 64:27]
  wire  _T_891; // @[Shift.scala 66:70]
  wire [26:0] _T_893; // @[Shift.scala 64:52]
  wire [27:0] _T_894; // @[Cat.scala 29:58]
  wire [27:0] _T_895; // @[Shift.scala 64:27]
  wire [27:0] _T_896; // @[Shift.scala 16:10]
  wire [2:0] _T_897; // @[convert.scala 23:34]
  wire [24:0] decC_fraction; // @[convert.scala 24:34]
  wire  _T_899; // @[convert.scala 25:26]
  wire [4:0] _T_901; // @[convert.scala 25:42]
  wire [2:0] _T_904; // @[convert.scala 26:67]
  wire [2:0] _T_905; // @[convert.scala 26:51]
  wire [8:0] _T_906; // @[Cat.scala 29:58]
  wire [29:0] _T_908; // @[convert.scala 29:56]
  wire  _T_909; // @[convert.scala 29:60]
  wire  _T_910; // @[convert.scala 29:41]
  wire  decC_isNaR; // @[convert.scala 29:39]
  wire  _T_913; // @[convert.scala 30:19]
  wire  decC_isZero; // @[convert.scala 30:41]
  wire [8:0] decC_scale; // @[convert.scala 32:24]
  wire  _T_921; // @[PositFMA.scala 58:30]
  wire  outIsNaR; // @[PositFMA.scala 58:44]
  wire  _T_922; // @[PositFMA.scala 59:34]
  wire  _T_923; // @[PositFMA.scala 59:47]
  wire  _T_924; // @[PositFMA.scala 59:45]
  wire [26:0] _T_926; // @[Cat.scala 29:58]
  wire [26:0] sigA; // @[PositFMA.scala 59:76]
  wire  _T_927; // @[PositFMA.scala 60:34]
  wire  _T_928; // @[PositFMA.scala 60:47]
  wire  _T_929; // @[PositFMA.scala 60:45]
  wire [26:0] _T_931; // @[Cat.scala 29:58]
  wire [26:0] sigB; // @[PositFMA.scala 60:76]
  wire [53:0] _T_932; // @[PositFMA.scala 61:25]
  wire [53:0] sigP; // @[PositFMA.scala 61:33]
  wire [1:0] head2; // @[PositFMA.scala 62:28]
  wire  _T_933; // @[PositFMA.scala 63:31]
  wire  _T_934; // @[PositFMA.scala 63:25]
  wire  _T_935; // @[PositFMA.scala 63:42]
  wire  addTwo; // @[PositFMA.scala 63:35]
  wire  _T_936; // @[PositFMA.scala 65:23]
  wire  _T_937; // @[PositFMA.scala 65:49]
  wire  addOne; // @[PositFMA.scala 65:43]
  wire [1:0] _T_938; // @[Cat.scala 29:58]
  wire [2:0] expBias; // @[PositFMA.scala 66:39]
  wire  mulSign; // @[PositFMA.scala 67:28]
  wire [9:0] _T_939; // @[PositFMA.scala 69:30]
  wire [9:0] _GEN_12; // @[PositFMA.scala 69:44]
  wire [9:0] _T_941; // @[PositFMA.scala 69:44]
  wire [9:0] mulScale; // @[PositFMA.scala 69:44]
  wire [51:0] _T_942; // @[PositFMA.scala 72:29]
  wire [50:0] _T_943; // @[PositFMA.scala 73:29]
  wire [51:0] _T_944; // @[PositFMA.scala 73:48]
  wire [51:0] mulSigTmp; // @[PositFMA.scala 70:22]
  wire  _T_946; // @[PositFMA.scala 77:39]
  wire  _T_947; // @[PositFMA.scala 77:43]
  wire [50:0] _T_948; // @[PositFMA.scala 78:39]
  wire [52:0] mulSig; // @[Cat.scala 29:58]
  reg  outIsNaR_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg [52:0] mulSig_phase2; // @[Reg.scala 15:16]
  reg [63:0] _RAND_1;
  reg [24:0] addFrac_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [9:0] mulScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [8:0] addScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  addSign_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  addZero_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  inValid_phase2; // @[Valid.scala 117:22]
  reg [31:0] _RAND_7;
  wire  _T_974; // @[PositFMA.scala 107:29]
  wire  _T_975; // @[PositFMA.scala 107:47]
  wire  _T_976; // @[PositFMA.scala 107:45]
  wire [52:0] extAddSig; // @[Cat.scala 29:58]
  wire [9:0] _GEN_13; // @[PositFMA.scala 111:39]
  wire  mulGreater; // @[PositFMA.scala 111:39]
  wire [9:0] greaterScale; // @[PositFMA.scala 112:26]
  wire [9:0] smallerScale; // @[PositFMA.scala 113:26]
  wire [9:0] _T_980; // @[PositFMA.scala 114:36]
  wire [9:0] scaleDiff; // @[PositFMA.scala 114:36]
  wire [52:0] greaterSig; // @[PositFMA.scala 115:26]
  wire [52:0] smallerSigTmp; // @[PositFMA.scala 116:26]
  wire [9:0] _T_981; // @[PositFMA.scala 117:69]
  wire  _T_982; // @[Shift.scala 39:24]
  wire [5:0] _T_983; // @[Shift.scala 40:44]
  wire [20:0] _T_984; // @[Shift.scala 90:30]
  wire [31:0] _T_985; // @[Shift.scala 90:48]
  wire  _T_986; // @[Shift.scala 90:57]
  wire [20:0] _GEN_14; // @[Shift.scala 90:39]
  wire [20:0] _T_987; // @[Shift.scala 90:39]
  wire  _T_988; // @[Shift.scala 12:21]
  wire  _T_989; // @[Shift.scala 12:21]
  wire [31:0] _T_991; // @[Bitwise.scala 71:12]
  wire [52:0] _T_992; // @[Cat.scala 29:58]
  wire [52:0] _T_993; // @[Shift.scala 91:22]
  wire [4:0] _T_994; // @[Shift.scala 92:77]
  wire [36:0] _T_995; // @[Shift.scala 90:30]
  wire [15:0] _T_996; // @[Shift.scala 90:48]
  wire  _T_997; // @[Shift.scala 90:57]
  wire [36:0] _GEN_15; // @[Shift.scala 90:39]
  wire [36:0] _T_998; // @[Shift.scala 90:39]
  wire  _T_999; // @[Shift.scala 12:21]
  wire  _T_1000; // @[Shift.scala 12:21]
  wire [15:0] _T_1002; // @[Bitwise.scala 71:12]
  wire [52:0] _T_1003; // @[Cat.scala 29:58]
  wire [52:0] _T_1004; // @[Shift.scala 91:22]
  wire [3:0] _T_1005; // @[Shift.scala 92:77]
  wire [44:0] _T_1006; // @[Shift.scala 90:30]
  wire [7:0] _T_1007; // @[Shift.scala 90:48]
  wire  _T_1008; // @[Shift.scala 90:57]
  wire [44:0] _GEN_16; // @[Shift.scala 90:39]
  wire [44:0] _T_1009; // @[Shift.scala 90:39]
  wire  _T_1010; // @[Shift.scala 12:21]
  wire  _T_1011; // @[Shift.scala 12:21]
  wire [7:0] _T_1013; // @[Bitwise.scala 71:12]
  wire [52:0] _T_1014; // @[Cat.scala 29:58]
  wire [52:0] _T_1015; // @[Shift.scala 91:22]
  wire [2:0] _T_1016; // @[Shift.scala 92:77]
  wire [48:0] _T_1017; // @[Shift.scala 90:30]
  wire [3:0] _T_1018; // @[Shift.scala 90:48]
  wire  _T_1019; // @[Shift.scala 90:57]
  wire [48:0] _GEN_17; // @[Shift.scala 90:39]
  wire [48:0] _T_1020; // @[Shift.scala 90:39]
  wire  _T_1021; // @[Shift.scala 12:21]
  wire  _T_1022; // @[Shift.scala 12:21]
  wire [3:0] _T_1024; // @[Bitwise.scala 71:12]
  wire [52:0] _T_1025; // @[Cat.scala 29:58]
  wire [52:0] _T_1026; // @[Shift.scala 91:22]
  wire [1:0] _T_1027; // @[Shift.scala 92:77]
  wire [50:0] _T_1028; // @[Shift.scala 90:30]
  wire [1:0] _T_1029; // @[Shift.scala 90:48]
  wire  _T_1030; // @[Shift.scala 90:57]
  wire [50:0] _GEN_18; // @[Shift.scala 90:39]
  wire [50:0] _T_1031; // @[Shift.scala 90:39]
  wire  _T_1032; // @[Shift.scala 12:21]
  wire  _T_1033; // @[Shift.scala 12:21]
  wire [1:0] _T_1035; // @[Bitwise.scala 71:12]
  wire [52:0] _T_1036; // @[Cat.scala 29:58]
  wire [52:0] _T_1037; // @[Shift.scala 91:22]
  wire  _T_1038; // @[Shift.scala 92:77]
  wire [51:0] _T_1039; // @[Shift.scala 90:30]
  wire  _T_1040; // @[Shift.scala 90:48]
  wire [51:0] _GEN_19; // @[Shift.scala 90:39]
  wire [51:0] _T_1042; // @[Shift.scala 90:39]
  wire  _T_1044; // @[Shift.scala 12:21]
  wire [52:0] _T_1045; // @[Cat.scala 29:58]
  wire [52:0] _T_1046; // @[Shift.scala 91:22]
  wire [52:0] _T_1049; // @[Bitwise.scala 71:12]
  wire [52:0] smallerSig; // @[Shift.scala 39:10]
  wire [53:0] rawSumSig; // @[PositFMA.scala 118:34]
  wire  _T_1050; // @[PositFMA.scala 119:42]
  wire  _T_1051; // @[PositFMA.scala 119:46]
  wire  _T_1052; // @[PositFMA.scala 119:79]
  wire  sumSign; // @[PositFMA.scala 119:63]
  wire [52:0] _T_1054; // @[PositFMA.scala 120:50]
  wire [53:0] signSumSig; // @[Cat.scala 29:58]
  wire [52:0] _T_1055; // @[PositFMA.scala 124:33]
  wire [52:0] _T_1056; // @[PositFMA.scala 124:68]
  wire [52:0] sumXor; // @[PositFMA.scala 124:51]
  wire [31:0] _T_1057; // @[LZD.scala 43:32]
  wire [15:0] _T_1058; // @[LZD.scala 43:32]
  wire [7:0] _T_1059; // @[LZD.scala 43:32]
  wire [3:0] _T_1060; // @[LZD.scala 43:32]
  wire [1:0] _T_1061; // @[LZD.scala 43:32]
  wire  _T_1062; // @[LZD.scala 39:14]
  wire  _T_1063; // @[LZD.scala 39:21]
  wire  _T_1064; // @[LZD.scala 39:30]
  wire  _T_1065; // @[LZD.scala 39:27]
  wire  _T_1066; // @[LZD.scala 39:25]
  wire [1:0] _T_1067; // @[Cat.scala 29:58]
  wire [1:0] _T_1068; // @[LZD.scala 44:32]
  wire  _T_1069; // @[LZD.scala 39:14]
  wire  _T_1070; // @[LZD.scala 39:21]
  wire  _T_1071; // @[LZD.scala 39:30]
  wire  _T_1072; // @[LZD.scala 39:27]
  wire  _T_1073; // @[LZD.scala 39:25]
  wire [1:0] _T_1074; // @[Cat.scala 29:58]
  wire  _T_1075; // @[Shift.scala 12:21]
  wire  _T_1076; // @[Shift.scala 12:21]
  wire  _T_1077; // @[LZD.scala 49:16]
  wire  _T_1078; // @[LZD.scala 49:27]
  wire  _T_1079; // @[LZD.scala 49:25]
  wire  _T_1080; // @[LZD.scala 49:47]
  wire  _T_1081; // @[LZD.scala 49:59]
  wire  _T_1082; // @[LZD.scala 49:35]
  wire [2:0] _T_1084; // @[Cat.scala 29:58]
  wire [3:0] _T_1085; // @[LZD.scala 44:32]
  wire [1:0] _T_1086; // @[LZD.scala 43:32]
  wire  _T_1087; // @[LZD.scala 39:14]
  wire  _T_1088; // @[LZD.scala 39:21]
  wire  _T_1089; // @[LZD.scala 39:30]
  wire  _T_1090; // @[LZD.scala 39:27]
  wire  _T_1091; // @[LZD.scala 39:25]
  wire [1:0] _T_1092; // @[Cat.scala 29:58]
  wire [1:0] _T_1093; // @[LZD.scala 44:32]
  wire  _T_1094; // @[LZD.scala 39:14]
  wire  _T_1095; // @[LZD.scala 39:21]
  wire  _T_1096; // @[LZD.scala 39:30]
  wire  _T_1097; // @[LZD.scala 39:27]
  wire  _T_1098; // @[LZD.scala 39:25]
  wire [1:0] _T_1099; // @[Cat.scala 29:58]
  wire  _T_1100; // @[Shift.scala 12:21]
  wire  _T_1101; // @[Shift.scala 12:21]
  wire  _T_1102; // @[LZD.scala 49:16]
  wire  _T_1103; // @[LZD.scala 49:27]
  wire  _T_1104; // @[LZD.scala 49:25]
  wire  _T_1105; // @[LZD.scala 49:47]
  wire  _T_1106; // @[LZD.scala 49:59]
  wire  _T_1107; // @[LZD.scala 49:35]
  wire [2:0] _T_1109; // @[Cat.scala 29:58]
  wire  _T_1110; // @[Shift.scala 12:21]
  wire  _T_1111; // @[Shift.scala 12:21]
  wire  _T_1112; // @[LZD.scala 49:16]
  wire  _T_1113; // @[LZD.scala 49:27]
  wire  _T_1114; // @[LZD.scala 49:25]
  wire [1:0] _T_1115; // @[LZD.scala 49:47]
  wire [1:0] _T_1116; // @[LZD.scala 49:59]
  wire [1:0] _T_1117; // @[LZD.scala 49:35]
  wire [3:0] _T_1119; // @[Cat.scala 29:58]
  wire [7:0] _T_1120; // @[LZD.scala 44:32]
  wire [3:0] _T_1121; // @[LZD.scala 43:32]
  wire [1:0] _T_1122; // @[LZD.scala 43:32]
  wire  _T_1123; // @[LZD.scala 39:14]
  wire  _T_1124; // @[LZD.scala 39:21]
  wire  _T_1125; // @[LZD.scala 39:30]
  wire  _T_1126; // @[LZD.scala 39:27]
  wire  _T_1127; // @[LZD.scala 39:25]
  wire [1:0] _T_1128; // @[Cat.scala 29:58]
  wire [1:0] _T_1129; // @[LZD.scala 44:32]
  wire  _T_1130; // @[LZD.scala 39:14]
  wire  _T_1131; // @[LZD.scala 39:21]
  wire  _T_1132; // @[LZD.scala 39:30]
  wire  _T_1133; // @[LZD.scala 39:27]
  wire  _T_1134; // @[LZD.scala 39:25]
  wire [1:0] _T_1135; // @[Cat.scala 29:58]
  wire  _T_1136; // @[Shift.scala 12:21]
  wire  _T_1137; // @[Shift.scala 12:21]
  wire  _T_1138; // @[LZD.scala 49:16]
  wire  _T_1139; // @[LZD.scala 49:27]
  wire  _T_1140; // @[LZD.scala 49:25]
  wire  _T_1141; // @[LZD.scala 49:47]
  wire  _T_1142; // @[LZD.scala 49:59]
  wire  _T_1143; // @[LZD.scala 49:35]
  wire [2:0] _T_1145; // @[Cat.scala 29:58]
  wire [3:0] _T_1146; // @[LZD.scala 44:32]
  wire [1:0] _T_1147; // @[LZD.scala 43:32]
  wire  _T_1148; // @[LZD.scala 39:14]
  wire  _T_1149; // @[LZD.scala 39:21]
  wire  _T_1150; // @[LZD.scala 39:30]
  wire  _T_1151; // @[LZD.scala 39:27]
  wire  _T_1152; // @[LZD.scala 39:25]
  wire [1:0] _T_1153; // @[Cat.scala 29:58]
  wire [1:0] _T_1154; // @[LZD.scala 44:32]
  wire  _T_1155; // @[LZD.scala 39:14]
  wire  _T_1156; // @[LZD.scala 39:21]
  wire  _T_1157; // @[LZD.scala 39:30]
  wire  _T_1158; // @[LZD.scala 39:27]
  wire  _T_1159; // @[LZD.scala 39:25]
  wire [1:0] _T_1160; // @[Cat.scala 29:58]
  wire  _T_1161; // @[Shift.scala 12:21]
  wire  _T_1162; // @[Shift.scala 12:21]
  wire  _T_1163; // @[LZD.scala 49:16]
  wire  _T_1164; // @[LZD.scala 49:27]
  wire  _T_1165; // @[LZD.scala 49:25]
  wire  _T_1166; // @[LZD.scala 49:47]
  wire  _T_1167; // @[LZD.scala 49:59]
  wire  _T_1168; // @[LZD.scala 49:35]
  wire [2:0] _T_1170; // @[Cat.scala 29:58]
  wire  _T_1171; // @[Shift.scala 12:21]
  wire  _T_1172; // @[Shift.scala 12:21]
  wire  _T_1173; // @[LZD.scala 49:16]
  wire  _T_1174; // @[LZD.scala 49:27]
  wire  _T_1175; // @[LZD.scala 49:25]
  wire [1:0] _T_1176; // @[LZD.scala 49:47]
  wire [1:0] _T_1177; // @[LZD.scala 49:59]
  wire [1:0] _T_1178; // @[LZD.scala 49:35]
  wire [3:0] _T_1180; // @[Cat.scala 29:58]
  wire  _T_1181; // @[Shift.scala 12:21]
  wire  _T_1182; // @[Shift.scala 12:21]
  wire  _T_1183; // @[LZD.scala 49:16]
  wire  _T_1184; // @[LZD.scala 49:27]
  wire  _T_1185; // @[LZD.scala 49:25]
  wire [2:0] _T_1186; // @[LZD.scala 49:47]
  wire [2:0] _T_1187; // @[LZD.scala 49:59]
  wire [2:0] _T_1188; // @[LZD.scala 49:35]
  wire [4:0] _T_1190; // @[Cat.scala 29:58]
  wire [15:0] _T_1191; // @[LZD.scala 44:32]
  wire [7:0] _T_1192; // @[LZD.scala 43:32]
  wire [3:0] _T_1193; // @[LZD.scala 43:32]
  wire [1:0] _T_1194; // @[LZD.scala 43:32]
  wire  _T_1195; // @[LZD.scala 39:14]
  wire  _T_1196; // @[LZD.scala 39:21]
  wire  _T_1197; // @[LZD.scala 39:30]
  wire  _T_1198; // @[LZD.scala 39:27]
  wire  _T_1199; // @[LZD.scala 39:25]
  wire [1:0] _T_1200; // @[Cat.scala 29:58]
  wire [1:0] _T_1201; // @[LZD.scala 44:32]
  wire  _T_1202; // @[LZD.scala 39:14]
  wire  _T_1203; // @[LZD.scala 39:21]
  wire  _T_1204; // @[LZD.scala 39:30]
  wire  _T_1205; // @[LZD.scala 39:27]
  wire  _T_1206; // @[LZD.scala 39:25]
  wire [1:0] _T_1207; // @[Cat.scala 29:58]
  wire  _T_1208; // @[Shift.scala 12:21]
  wire  _T_1209; // @[Shift.scala 12:21]
  wire  _T_1210; // @[LZD.scala 49:16]
  wire  _T_1211; // @[LZD.scala 49:27]
  wire  _T_1212; // @[LZD.scala 49:25]
  wire  _T_1213; // @[LZD.scala 49:47]
  wire  _T_1214; // @[LZD.scala 49:59]
  wire  _T_1215; // @[LZD.scala 49:35]
  wire [2:0] _T_1217; // @[Cat.scala 29:58]
  wire [3:0] _T_1218; // @[LZD.scala 44:32]
  wire [1:0] _T_1219; // @[LZD.scala 43:32]
  wire  _T_1220; // @[LZD.scala 39:14]
  wire  _T_1221; // @[LZD.scala 39:21]
  wire  _T_1222; // @[LZD.scala 39:30]
  wire  _T_1223; // @[LZD.scala 39:27]
  wire  _T_1224; // @[LZD.scala 39:25]
  wire [1:0] _T_1225; // @[Cat.scala 29:58]
  wire [1:0] _T_1226; // @[LZD.scala 44:32]
  wire  _T_1227; // @[LZD.scala 39:14]
  wire  _T_1228; // @[LZD.scala 39:21]
  wire  _T_1229; // @[LZD.scala 39:30]
  wire  _T_1230; // @[LZD.scala 39:27]
  wire  _T_1231; // @[LZD.scala 39:25]
  wire [1:0] _T_1232; // @[Cat.scala 29:58]
  wire  _T_1233; // @[Shift.scala 12:21]
  wire  _T_1234; // @[Shift.scala 12:21]
  wire  _T_1235; // @[LZD.scala 49:16]
  wire  _T_1236; // @[LZD.scala 49:27]
  wire  _T_1237; // @[LZD.scala 49:25]
  wire  _T_1238; // @[LZD.scala 49:47]
  wire  _T_1239; // @[LZD.scala 49:59]
  wire  _T_1240; // @[LZD.scala 49:35]
  wire [2:0] _T_1242; // @[Cat.scala 29:58]
  wire  _T_1243; // @[Shift.scala 12:21]
  wire  _T_1244; // @[Shift.scala 12:21]
  wire  _T_1245; // @[LZD.scala 49:16]
  wire  _T_1246; // @[LZD.scala 49:27]
  wire  _T_1247; // @[LZD.scala 49:25]
  wire [1:0] _T_1248; // @[LZD.scala 49:47]
  wire [1:0] _T_1249; // @[LZD.scala 49:59]
  wire [1:0] _T_1250; // @[LZD.scala 49:35]
  wire [3:0] _T_1252; // @[Cat.scala 29:58]
  wire [7:0] _T_1253; // @[LZD.scala 44:32]
  wire [3:0] _T_1254; // @[LZD.scala 43:32]
  wire [1:0] _T_1255; // @[LZD.scala 43:32]
  wire  _T_1256; // @[LZD.scala 39:14]
  wire  _T_1257; // @[LZD.scala 39:21]
  wire  _T_1258; // @[LZD.scala 39:30]
  wire  _T_1259; // @[LZD.scala 39:27]
  wire  _T_1260; // @[LZD.scala 39:25]
  wire [1:0] _T_1261; // @[Cat.scala 29:58]
  wire [1:0] _T_1262; // @[LZD.scala 44:32]
  wire  _T_1263; // @[LZD.scala 39:14]
  wire  _T_1264; // @[LZD.scala 39:21]
  wire  _T_1265; // @[LZD.scala 39:30]
  wire  _T_1266; // @[LZD.scala 39:27]
  wire  _T_1267; // @[LZD.scala 39:25]
  wire [1:0] _T_1268; // @[Cat.scala 29:58]
  wire  _T_1269; // @[Shift.scala 12:21]
  wire  _T_1270; // @[Shift.scala 12:21]
  wire  _T_1271; // @[LZD.scala 49:16]
  wire  _T_1272; // @[LZD.scala 49:27]
  wire  _T_1273; // @[LZD.scala 49:25]
  wire  _T_1274; // @[LZD.scala 49:47]
  wire  _T_1275; // @[LZD.scala 49:59]
  wire  _T_1276; // @[LZD.scala 49:35]
  wire [2:0] _T_1278; // @[Cat.scala 29:58]
  wire [3:0] _T_1279; // @[LZD.scala 44:32]
  wire [1:0] _T_1280; // @[LZD.scala 43:32]
  wire  _T_1281; // @[LZD.scala 39:14]
  wire  _T_1282; // @[LZD.scala 39:21]
  wire  _T_1283; // @[LZD.scala 39:30]
  wire  _T_1284; // @[LZD.scala 39:27]
  wire  _T_1285; // @[LZD.scala 39:25]
  wire [1:0] _T_1286; // @[Cat.scala 29:58]
  wire [1:0] _T_1287; // @[LZD.scala 44:32]
  wire  _T_1288; // @[LZD.scala 39:14]
  wire  _T_1289; // @[LZD.scala 39:21]
  wire  _T_1290; // @[LZD.scala 39:30]
  wire  _T_1291; // @[LZD.scala 39:27]
  wire  _T_1292; // @[LZD.scala 39:25]
  wire [1:0] _T_1293; // @[Cat.scala 29:58]
  wire  _T_1294; // @[Shift.scala 12:21]
  wire  _T_1295; // @[Shift.scala 12:21]
  wire  _T_1296; // @[LZD.scala 49:16]
  wire  _T_1297; // @[LZD.scala 49:27]
  wire  _T_1298; // @[LZD.scala 49:25]
  wire  _T_1299; // @[LZD.scala 49:47]
  wire  _T_1300; // @[LZD.scala 49:59]
  wire  _T_1301; // @[LZD.scala 49:35]
  wire [2:0] _T_1303; // @[Cat.scala 29:58]
  wire  _T_1304; // @[Shift.scala 12:21]
  wire  _T_1305; // @[Shift.scala 12:21]
  wire  _T_1306; // @[LZD.scala 49:16]
  wire  _T_1307; // @[LZD.scala 49:27]
  wire  _T_1308; // @[LZD.scala 49:25]
  wire [1:0] _T_1309; // @[LZD.scala 49:47]
  wire [1:0] _T_1310; // @[LZD.scala 49:59]
  wire [1:0] _T_1311; // @[LZD.scala 49:35]
  wire [3:0] _T_1313; // @[Cat.scala 29:58]
  wire  _T_1314; // @[Shift.scala 12:21]
  wire  _T_1315; // @[Shift.scala 12:21]
  wire  _T_1316; // @[LZD.scala 49:16]
  wire  _T_1317; // @[LZD.scala 49:27]
  wire  _T_1318; // @[LZD.scala 49:25]
  wire [2:0] _T_1319; // @[LZD.scala 49:47]
  wire [2:0] _T_1320; // @[LZD.scala 49:59]
  wire [2:0] _T_1321; // @[LZD.scala 49:35]
  wire [4:0] _T_1323; // @[Cat.scala 29:58]
  wire  _T_1324; // @[Shift.scala 12:21]
  wire  _T_1325; // @[Shift.scala 12:21]
  wire  _T_1326; // @[LZD.scala 49:16]
  wire  _T_1327; // @[LZD.scala 49:27]
  wire  _T_1328; // @[LZD.scala 49:25]
  wire [3:0] _T_1329; // @[LZD.scala 49:47]
  wire [3:0] _T_1330; // @[LZD.scala 49:59]
  wire [3:0] _T_1331; // @[LZD.scala 49:35]
  wire [5:0] _T_1333; // @[Cat.scala 29:58]
  wire [20:0] _T_1334; // @[LZD.scala 44:32]
  wire [15:0] _T_1335; // @[LZD.scala 43:32]
  wire [7:0] _T_1336; // @[LZD.scala 43:32]
  wire [3:0] _T_1337; // @[LZD.scala 43:32]
  wire [1:0] _T_1338; // @[LZD.scala 43:32]
  wire  _T_1339; // @[LZD.scala 39:14]
  wire  _T_1340; // @[LZD.scala 39:21]
  wire  _T_1341; // @[LZD.scala 39:30]
  wire  _T_1342; // @[LZD.scala 39:27]
  wire  _T_1343; // @[LZD.scala 39:25]
  wire [1:0] _T_1344; // @[Cat.scala 29:58]
  wire [1:0] _T_1345; // @[LZD.scala 44:32]
  wire  _T_1346; // @[LZD.scala 39:14]
  wire  _T_1347; // @[LZD.scala 39:21]
  wire  _T_1348; // @[LZD.scala 39:30]
  wire  _T_1349; // @[LZD.scala 39:27]
  wire  _T_1350; // @[LZD.scala 39:25]
  wire [1:0] _T_1351; // @[Cat.scala 29:58]
  wire  _T_1352; // @[Shift.scala 12:21]
  wire  _T_1353; // @[Shift.scala 12:21]
  wire  _T_1354; // @[LZD.scala 49:16]
  wire  _T_1355; // @[LZD.scala 49:27]
  wire  _T_1356; // @[LZD.scala 49:25]
  wire  _T_1357; // @[LZD.scala 49:47]
  wire  _T_1358; // @[LZD.scala 49:59]
  wire  _T_1359; // @[LZD.scala 49:35]
  wire [2:0] _T_1361; // @[Cat.scala 29:58]
  wire [3:0] _T_1362; // @[LZD.scala 44:32]
  wire [1:0] _T_1363; // @[LZD.scala 43:32]
  wire  _T_1364; // @[LZD.scala 39:14]
  wire  _T_1365; // @[LZD.scala 39:21]
  wire  _T_1366; // @[LZD.scala 39:30]
  wire  _T_1367; // @[LZD.scala 39:27]
  wire  _T_1368; // @[LZD.scala 39:25]
  wire [1:0] _T_1369; // @[Cat.scala 29:58]
  wire [1:0] _T_1370; // @[LZD.scala 44:32]
  wire  _T_1371; // @[LZD.scala 39:14]
  wire  _T_1372; // @[LZD.scala 39:21]
  wire  _T_1373; // @[LZD.scala 39:30]
  wire  _T_1374; // @[LZD.scala 39:27]
  wire  _T_1375; // @[LZD.scala 39:25]
  wire [1:0] _T_1376; // @[Cat.scala 29:58]
  wire  _T_1377; // @[Shift.scala 12:21]
  wire  _T_1378; // @[Shift.scala 12:21]
  wire  _T_1379; // @[LZD.scala 49:16]
  wire  _T_1380; // @[LZD.scala 49:27]
  wire  _T_1381; // @[LZD.scala 49:25]
  wire  _T_1382; // @[LZD.scala 49:47]
  wire  _T_1383; // @[LZD.scala 49:59]
  wire  _T_1384; // @[LZD.scala 49:35]
  wire [2:0] _T_1386; // @[Cat.scala 29:58]
  wire  _T_1387; // @[Shift.scala 12:21]
  wire  _T_1388; // @[Shift.scala 12:21]
  wire  _T_1389; // @[LZD.scala 49:16]
  wire  _T_1390; // @[LZD.scala 49:27]
  wire  _T_1391; // @[LZD.scala 49:25]
  wire [1:0] _T_1392; // @[LZD.scala 49:47]
  wire [1:0] _T_1393; // @[LZD.scala 49:59]
  wire [1:0] _T_1394; // @[LZD.scala 49:35]
  wire [3:0] _T_1396; // @[Cat.scala 29:58]
  wire [7:0] _T_1397; // @[LZD.scala 44:32]
  wire [3:0] _T_1398; // @[LZD.scala 43:32]
  wire [1:0] _T_1399; // @[LZD.scala 43:32]
  wire  _T_1400; // @[LZD.scala 39:14]
  wire  _T_1401; // @[LZD.scala 39:21]
  wire  _T_1402; // @[LZD.scala 39:30]
  wire  _T_1403; // @[LZD.scala 39:27]
  wire  _T_1404; // @[LZD.scala 39:25]
  wire [1:0] _T_1405; // @[Cat.scala 29:58]
  wire [1:0] _T_1406; // @[LZD.scala 44:32]
  wire  _T_1407; // @[LZD.scala 39:14]
  wire  _T_1408; // @[LZD.scala 39:21]
  wire  _T_1409; // @[LZD.scala 39:30]
  wire  _T_1410; // @[LZD.scala 39:27]
  wire  _T_1411; // @[LZD.scala 39:25]
  wire [1:0] _T_1412; // @[Cat.scala 29:58]
  wire  _T_1413; // @[Shift.scala 12:21]
  wire  _T_1414; // @[Shift.scala 12:21]
  wire  _T_1415; // @[LZD.scala 49:16]
  wire  _T_1416; // @[LZD.scala 49:27]
  wire  _T_1417; // @[LZD.scala 49:25]
  wire  _T_1418; // @[LZD.scala 49:47]
  wire  _T_1419; // @[LZD.scala 49:59]
  wire  _T_1420; // @[LZD.scala 49:35]
  wire [2:0] _T_1422; // @[Cat.scala 29:58]
  wire [3:0] _T_1423; // @[LZD.scala 44:32]
  wire [1:0] _T_1424; // @[LZD.scala 43:32]
  wire  _T_1425; // @[LZD.scala 39:14]
  wire  _T_1426; // @[LZD.scala 39:21]
  wire  _T_1427; // @[LZD.scala 39:30]
  wire  _T_1428; // @[LZD.scala 39:27]
  wire  _T_1429; // @[LZD.scala 39:25]
  wire [1:0] _T_1430; // @[Cat.scala 29:58]
  wire [1:0] _T_1431; // @[LZD.scala 44:32]
  wire  _T_1432; // @[LZD.scala 39:14]
  wire  _T_1433; // @[LZD.scala 39:21]
  wire  _T_1434; // @[LZD.scala 39:30]
  wire  _T_1435; // @[LZD.scala 39:27]
  wire  _T_1436; // @[LZD.scala 39:25]
  wire [1:0] _T_1437; // @[Cat.scala 29:58]
  wire  _T_1438; // @[Shift.scala 12:21]
  wire  _T_1439; // @[Shift.scala 12:21]
  wire  _T_1440; // @[LZD.scala 49:16]
  wire  _T_1441; // @[LZD.scala 49:27]
  wire  _T_1442; // @[LZD.scala 49:25]
  wire  _T_1443; // @[LZD.scala 49:47]
  wire  _T_1444; // @[LZD.scala 49:59]
  wire  _T_1445; // @[LZD.scala 49:35]
  wire [2:0] _T_1447; // @[Cat.scala 29:58]
  wire  _T_1448; // @[Shift.scala 12:21]
  wire  _T_1449; // @[Shift.scala 12:21]
  wire  _T_1450; // @[LZD.scala 49:16]
  wire  _T_1451; // @[LZD.scala 49:27]
  wire  _T_1452; // @[LZD.scala 49:25]
  wire [1:0] _T_1453; // @[LZD.scala 49:47]
  wire [1:0] _T_1454; // @[LZD.scala 49:59]
  wire [1:0] _T_1455; // @[LZD.scala 49:35]
  wire [3:0] _T_1457; // @[Cat.scala 29:58]
  wire  _T_1458; // @[Shift.scala 12:21]
  wire  _T_1459; // @[Shift.scala 12:21]
  wire  _T_1460; // @[LZD.scala 49:16]
  wire  _T_1461; // @[LZD.scala 49:27]
  wire  _T_1462; // @[LZD.scala 49:25]
  wire [2:0] _T_1463; // @[LZD.scala 49:47]
  wire [2:0] _T_1464; // @[LZD.scala 49:59]
  wire [2:0] _T_1465; // @[LZD.scala 49:35]
  wire [4:0] _T_1467; // @[Cat.scala 29:58]
  wire [4:0] _T_1468; // @[LZD.scala 44:32]
  wire [3:0] _T_1469; // @[LZD.scala 43:32]
  wire [1:0] _T_1470; // @[LZD.scala 43:32]
  wire  _T_1471; // @[LZD.scala 39:14]
  wire  _T_1472; // @[LZD.scala 39:21]
  wire  _T_1473; // @[LZD.scala 39:30]
  wire  _T_1474; // @[LZD.scala 39:27]
  wire  _T_1475; // @[LZD.scala 39:25]
  wire [1:0] _T_1476; // @[Cat.scala 29:58]
  wire [1:0] _T_1477; // @[LZD.scala 44:32]
  wire  _T_1478; // @[LZD.scala 39:14]
  wire  _T_1479; // @[LZD.scala 39:21]
  wire  _T_1480; // @[LZD.scala 39:30]
  wire  _T_1481; // @[LZD.scala 39:27]
  wire  _T_1482; // @[LZD.scala 39:25]
  wire [1:0] _T_1483; // @[Cat.scala 29:58]
  wire  _T_1484; // @[Shift.scala 12:21]
  wire  _T_1485; // @[Shift.scala 12:21]
  wire  _T_1486; // @[LZD.scala 49:16]
  wire  _T_1487; // @[LZD.scala 49:27]
  wire  _T_1488; // @[LZD.scala 49:25]
  wire  _T_1489; // @[LZD.scala 49:47]
  wire  _T_1490; // @[LZD.scala 49:59]
  wire  _T_1491; // @[LZD.scala 49:35]
  wire [2:0] _T_1493; // @[Cat.scala 29:58]
  wire  _T_1494; // @[LZD.scala 44:32]
  wire  _T_1496; // @[Shift.scala 12:21]
  wire [1:0] _T_1498; // @[Cat.scala 29:58]
  wire [1:0] _T_1499; // @[LZD.scala 55:32]
  wire [1:0] _T_1500; // @[LZD.scala 55:20]
  wire  _T_1502; // @[Shift.scala 12:21]
  wire [3:0] _T_1504; // @[Cat.scala 29:58]
  wire [3:0] _T_1505; // @[LZD.scala 55:32]
  wire [3:0] _T_1506; // @[LZD.scala 55:20]
  wire [4:0] _T_1507; // @[Cat.scala 29:58]
  wire  _T_1508; // @[Shift.scala 12:21]
  wire [4:0] _T_1510; // @[LZD.scala 55:32]
  wire [4:0] _T_1511; // @[LZD.scala 55:20]
  wire [5:0] sumLZD; // @[Cat.scala 29:58]
  wire [5:0] shiftValue; // @[PositFMA.scala 126:24]
  wire [51:0] _T_1512; // @[PositFMA.scala 127:38]
  wire  _T_1513; // @[Shift.scala 16:24]
  wire  _T_1515; // @[Shift.scala 12:21]
  wire [19:0] _T_1516; // @[Shift.scala 64:52]
  wire [51:0] _T_1518; // @[Cat.scala 29:58]
  wire [51:0] _T_1519; // @[Shift.scala 64:27]
  wire [4:0] _T_1520; // @[Shift.scala 66:70]
  wire  _T_1521; // @[Shift.scala 12:21]
  wire [35:0] _T_1522; // @[Shift.scala 64:52]
  wire [51:0] _T_1524; // @[Cat.scala 29:58]
  wire [51:0] _T_1525; // @[Shift.scala 64:27]
  wire [3:0] _T_1526; // @[Shift.scala 66:70]
  wire  _T_1527; // @[Shift.scala 12:21]
  wire [43:0] _T_1528; // @[Shift.scala 64:52]
  wire [51:0] _T_1530; // @[Cat.scala 29:58]
  wire [51:0] _T_1531; // @[Shift.scala 64:27]
  wire [2:0] _T_1532; // @[Shift.scala 66:70]
  wire  _T_1533; // @[Shift.scala 12:21]
  wire [47:0] _T_1534; // @[Shift.scala 64:52]
  wire [51:0] _T_1536; // @[Cat.scala 29:58]
  wire [51:0] _T_1537; // @[Shift.scala 64:27]
  wire [1:0] _T_1538; // @[Shift.scala 66:70]
  wire  _T_1539; // @[Shift.scala 12:21]
  wire [49:0] _T_1540; // @[Shift.scala 64:52]
  wire [51:0] _T_1542; // @[Cat.scala 29:58]
  wire [51:0] _T_1543; // @[Shift.scala 64:27]
  wire  _T_1544; // @[Shift.scala 66:70]
  wire [50:0] _T_1546; // @[Shift.scala 64:52]
  wire [51:0] _T_1547; // @[Cat.scala 29:58]
  wire [51:0] _T_1548; // @[Shift.scala 64:27]
  wire [51:0] normalFracTmp; // @[Shift.scala 16:10]
  wire [9:0] _T_1550; // @[PositFMA.scala 130:36]
  wire [9:0] _T_1551; // @[PositFMA.scala 130:36]
  wire [6:0] _T_1552; // @[Cat.scala 29:58]
  wire [6:0] _T_1553; // @[PositFMA.scala 130:61]
  wire [9:0] _GEN_20; // @[PositFMA.scala 130:42]
  wire [9:0] _T_1555; // @[PositFMA.scala 130:42]
  wire [9:0] sumScale; // @[PositFMA.scala 130:42]
  wire [24:0] sumFrac; // @[PositFMA.scala 131:41]
  wire [26:0] grsTmp; // @[PositFMA.scala 134:41]
  wire [1:0] _T_1556; // @[PositFMA.scala 137:40]
  wire [24:0] _T_1557; // @[PositFMA.scala 137:56]
  wire  _T_1558; // @[PositFMA.scala 137:60]
  wire  underflow; // @[PositFMA.scala 144:32]
  wire  overflow; // @[PositFMA.scala 145:32]
  wire  _T_1559; // @[PositFMA.scala 154:32]
  wire  decF_isZero; // @[PositFMA.scala 154:20]
  wire [9:0] _T_1561; // @[Mux.scala 87:16]
  wire [9:0] _T_1562; // @[Mux.scala 87:16]
  wire [8:0] _GEN_21; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  wire [8:0] decF_scale; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  wire [2:0] _T_1563; // @[convert.scala 46:61]
  wire [2:0] _T_1564; // @[convert.scala 46:52]
  wire [2:0] _T_1566; // @[convert.scala 46:42]
  wire [5:0] _T_1567; // @[convert.scala 48:34]
  wire  _T_1568; // @[convert.scala 49:36]
  wire [5:0] _T_1570; // @[convert.scala 50:36]
  wire [5:0] _T_1571; // @[convert.scala 50:36]
  wire [5:0] _T_1572; // @[convert.scala 50:28]
  wire  _T_1573; // @[convert.scala 51:31]
  wire  _T_1574; // @[convert.scala 52:43]
  wire [32:0] _T_1578; // @[Cat.scala 29:58]
  wire [5:0] _T_1579; // @[Shift.scala 39:17]
  wire  _T_1580; // @[Shift.scala 39:24]
  wire  _T_1582; // @[Shift.scala 90:30]
  wire [31:0] _T_1583; // @[Shift.scala 90:48]
  wire  _T_1584; // @[Shift.scala 90:57]
  wire  _T_1585; // @[Shift.scala 90:39]
  wire  _T_1586; // @[Shift.scala 12:21]
  wire  _T_1587; // @[Shift.scala 12:21]
  wire [31:0] _T_1589; // @[Bitwise.scala 71:12]
  wire [32:0] _T_1590; // @[Cat.scala 29:58]
  wire [32:0] _T_1591; // @[Shift.scala 91:22]
  wire [4:0] _T_1592; // @[Shift.scala 92:77]
  wire [16:0] _T_1593; // @[Shift.scala 90:30]
  wire [15:0] _T_1594; // @[Shift.scala 90:48]
  wire  _T_1595; // @[Shift.scala 90:57]
  wire [16:0] _GEN_22; // @[Shift.scala 90:39]
  wire [16:0] _T_1596; // @[Shift.scala 90:39]
  wire  _T_1597; // @[Shift.scala 12:21]
  wire  _T_1598; // @[Shift.scala 12:21]
  wire [15:0] _T_1600; // @[Bitwise.scala 71:12]
  wire [32:0] _T_1601; // @[Cat.scala 29:58]
  wire [32:0] _T_1602; // @[Shift.scala 91:22]
  wire [3:0] _T_1603; // @[Shift.scala 92:77]
  wire [24:0] _T_1604; // @[Shift.scala 90:30]
  wire [7:0] _T_1605; // @[Shift.scala 90:48]
  wire  _T_1606; // @[Shift.scala 90:57]
  wire [24:0] _GEN_23; // @[Shift.scala 90:39]
  wire [24:0] _T_1607; // @[Shift.scala 90:39]
  wire  _T_1608; // @[Shift.scala 12:21]
  wire  _T_1609; // @[Shift.scala 12:21]
  wire [7:0] _T_1611; // @[Bitwise.scala 71:12]
  wire [32:0] _T_1612; // @[Cat.scala 29:58]
  wire [32:0] _T_1613; // @[Shift.scala 91:22]
  wire [2:0] _T_1614; // @[Shift.scala 92:77]
  wire [28:0] _T_1615; // @[Shift.scala 90:30]
  wire [3:0] _T_1616; // @[Shift.scala 90:48]
  wire  _T_1617; // @[Shift.scala 90:57]
  wire [28:0] _GEN_24; // @[Shift.scala 90:39]
  wire [28:0] _T_1618; // @[Shift.scala 90:39]
  wire  _T_1619; // @[Shift.scala 12:21]
  wire  _T_1620; // @[Shift.scala 12:21]
  wire [3:0] _T_1622; // @[Bitwise.scala 71:12]
  wire [32:0] _T_1623; // @[Cat.scala 29:58]
  wire [32:0] _T_1624; // @[Shift.scala 91:22]
  wire [1:0] _T_1625; // @[Shift.scala 92:77]
  wire [30:0] _T_1626; // @[Shift.scala 90:30]
  wire [1:0] _T_1627; // @[Shift.scala 90:48]
  wire  _T_1628; // @[Shift.scala 90:57]
  wire [30:0] _GEN_25; // @[Shift.scala 90:39]
  wire [30:0] _T_1629; // @[Shift.scala 90:39]
  wire  _T_1630; // @[Shift.scala 12:21]
  wire  _T_1631; // @[Shift.scala 12:21]
  wire [1:0] _T_1633; // @[Bitwise.scala 71:12]
  wire [32:0] _T_1634; // @[Cat.scala 29:58]
  wire [32:0] _T_1635; // @[Shift.scala 91:22]
  wire  _T_1636; // @[Shift.scala 92:77]
  wire [31:0] _T_1637; // @[Shift.scala 90:30]
  wire  _T_1638; // @[Shift.scala 90:48]
  wire [31:0] _GEN_26; // @[Shift.scala 90:39]
  wire [31:0] _T_1640; // @[Shift.scala 90:39]
  wire  _T_1642; // @[Shift.scala 12:21]
  wire [32:0] _T_1643; // @[Cat.scala 29:58]
  wire [32:0] _T_1644; // @[Shift.scala 91:22]
  wire [32:0] _T_1647; // @[Bitwise.scala 71:12]
  wire [32:0] _T_1648; // @[Shift.scala 39:10]
  wire  _T_1649; // @[convert.scala 55:31]
  wire  _T_1650; // @[convert.scala 56:31]
  wire  _T_1651; // @[convert.scala 57:31]
  wire  _T_1652; // @[convert.scala 58:31]
  wire [29:0] _T_1653; // @[convert.scala 59:69]
  wire  _T_1654; // @[convert.scala 59:81]
  wire  _T_1655; // @[convert.scala 59:50]
  wire  _T_1657; // @[convert.scala 60:81]
  wire  _T_1658; // @[convert.scala 61:44]
  wire  _T_1659; // @[convert.scala 61:52]
  wire  _T_1660; // @[convert.scala 61:36]
  wire  _T_1661; // @[convert.scala 62:63]
  wire  _T_1662; // @[convert.scala 62:103]
  wire  _T_1663; // @[convert.scala 62:60]
  wire [29:0] _GEN_27; // @[convert.scala 63:56]
  wire [29:0] _T_1666; // @[convert.scala 63:56]
  wire [30:0] _T_1667; // @[Cat.scala 29:58]
  reg  _T_1671; // @[Valid.scala 117:22]
  reg [31:0] _RAND_8;
  reg [30:0] _T_1675; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  assign _T = io_fmaOp[1]; // @[PositFMA.scala 47:36]
  assign _T_2 = _T ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 71:12]
  assign _T_3 = _T_2 ^ io_A; // @[PositFMA.scala 47:41]
  assign _GEN_10 = {{30'd0}, _T}; // @[PositFMA.scala 47:49]
  assign realA = _T_3 + _GEN_10; // @[PositFMA.scala 47:49]
  assign _T_6 = io_fmaOp[0]; // @[PositFMA.scala 48:36]
  assign _T_8 = _T_6 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 71:12]
  assign _T_9 = _T_8 ^ io_C; // @[PositFMA.scala 48:41]
  assign _GEN_11 = {{30'd0}, _T_6}; // @[PositFMA.scala 48:49]
  assign realC = _T_9 + _GEN_11; // @[PositFMA.scala 48:49]
  assign _T_13 = realA[30]; // @[convert.scala 18:24]
  assign _T_14 = realA[29]; // @[convert.scala 18:40]
  assign _T_15 = _T_13 ^ _T_14; // @[convert.scala 18:36]
  assign _T_16 = realA[29:1]; // @[convert.scala 19:24]
  assign _T_17 = realA[28:0]; // @[convert.scala 19:43]
  assign _T_18 = _T_16 ^ _T_17; // @[convert.scala 19:39]
  assign _T_19 = _T_18[28:13]; // @[LZD.scala 43:32]
  assign _T_20 = _T_19[15:8]; // @[LZD.scala 43:32]
  assign _T_21 = _T_20[7:4]; // @[LZD.scala 43:32]
  assign _T_22 = _T_21[3:2]; // @[LZD.scala 43:32]
  assign _T_23 = _T_22 != 2'h0; // @[LZD.scala 39:14]
  assign _T_24 = _T_22[1]; // @[LZD.scala 39:21]
  assign _T_25 = _T_22[0]; // @[LZD.scala 39:30]
  assign _T_26 = ~ _T_25; // @[LZD.scala 39:27]
  assign _T_27 = _T_24 | _T_26; // @[LZD.scala 39:25]
  assign _T_28 = {_T_23,_T_27}; // @[Cat.scala 29:58]
  assign _T_29 = _T_21[1:0]; // @[LZD.scala 44:32]
  assign _T_30 = _T_29 != 2'h0; // @[LZD.scala 39:14]
  assign _T_31 = _T_29[1]; // @[LZD.scala 39:21]
  assign _T_32 = _T_29[0]; // @[LZD.scala 39:30]
  assign _T_33 = ~ _T_32; // @[LZD.scala 39:27]
  assign _T_34 = _T_31 | _T_33; // @[LZD.scala 39:25]
  assign _T_35 = {_T_30,_T_34}; // @[Cat.scala 29:58]
  assign _T_36 = _T_28[1]; // @[Shift.scala 12:21]
  assign _T_37 = _T_35[1]; // @[Shift.scala 12:21]
  assign _T_38 = _T_36 | _T_37; // @[LZD.scala 49:16]
  assign _T_39 = ~ _T_37; // @[LZD.scala 49:27]
  assign _T_40 = _T_36 | _T_39; // @[LZD.scala 49:25]
  assign _T_41 = _T_28[0:0]; // @[LZD.scala 49:47]
  assign _T_42 = _T_35[0:0]; // @[LZD.scala 49:59]
  assign _T_43 = _T_36 ? _T_41 : _T_42; // @[LZD.scala 49:35]
  assign _T_45 = {_T_38,_T_40,_T_43}; // @[Cat.scala 29:58]
  assign _T_46 = _T_20[3:0]; // @[LZD.scala 44:32]
  assign _T_47 = _T_46[3:2]; // @[LZD.scala 43:32]
  assign _T_48 = _T_47 != 2'h0; // @[LZD.scala 39:14]
  assign _T_49 = _T_47[1]; // @[LZD.scala 39:21]
  assign _T_50 = _T_47[0]; // @[LZD.scala 39:30]
  assign _T_51 = ~ _T_50; // @[LZD.scala 39:27]
  assign _T_52 = _T_49 | _T_51; // @[LZD.scala 39:25]
  assign _T_53 = {_T_48,_T_52}; // @[Cat.scala 29:58]
  assign _T_54 = _T_46[1:0]; // @[LZD.scala 44:32]
  assign _T_55 = _T_54 != 2'h0; // @[LZD.scala 39:14]
  assign _T_56 = _T_54[1]; // @[LZD.scala 39:21]
  assign _T_57 = _T_54[0]; // @[LZD.scala 39:30]
  assign _T_58 = ~ _T_57; // @[LZD.scala 39:27]
  assign _T_59 = _T_56 | _T_58; // @[LZD.scala 39:25]
  assign _T_60 = {_T_55,_T_59}; // @[Cat.scala 29:58]
  assign _T_61 = _T_53[1]; // @[Shift.scala 12:21]
  assign _T_62 = _T_60[1]; // @[Shift.scala 12:21]
  assign _T_63 = _T_61 | _T_62; // @[LZD.scala 49:16]
  assign _T_64 = ~ _T_62; // @[LZD.scala 49:27]
  assign _T_65 = _T_61 | _T_64; // @[LZD.scala 49:25]
  assign _T_66 = _T_53[0:0]; // @[LZD.scala 49:47]
  assign _T_67 = _T_60[0:0]; // @[LZD.scala 49:59]
  assign _T_68 = _T_61 ? _T_66 : _T_67; // @[LZD.scala 49:35]
  assign _T_70 = {_T_63,_T_65,_T_68}; // @[Cat.scala 29:58]
  assign _T_71 = _T_45[2]; // @[Shift.scala 12:21]
  assign _T_72 = _T_70[2]; // @[Shift.scala 12:21]
  assign _T_73 = _T_71 | _T_72; // @[LZD.scala 49:16]
  assign _T_74 = ~ _T_72; // @[LZD.scala 49:27]
  assign _T_75 = _T_71 | _T_74; // @[LZD.scala 49:25]
  assign _T_76 = _T_45[1:0]; // @[LZD.scala 49:47]
  assign _T_77 = _T_70[1:0]; // @[LZD.scala 49:59]
  assign _T_78 = _T_71 ? _T_76 : _T_77; // @[LZD.scala 49:35]
  assign _T_80 = {_T_73,_T_75,_T_78}; // @[Cat.scala 29:58]
  assign _T_81 = _T_19[7:0]; // @[LZD.scala 44:32]
  assign _T_82 = _T_81[7:4]; // @[LZD.scala 43:32]
  assign _T_83 = _T_82[3:2]; // @[LZD.scala 43:32]
  assign _T_84 = _T_83 != 2'h0; // @[LZD.scala 39:14]
  assign _T_85 = _T_83[1]; // @[LZD.scala 39:21]
  assign _T_86 = _T_83[0]; // @[LZD.scala 39:30]
  assign _T_87 = ~ _T_86; // @[LZD.scala 39:27]
  assign _T_88 = _T_85 | _T_87; // @[LZD.scala 39:25]
  assign _T_89 = {_T_84,_T_88}; // @[Cat.scala 29:58]
  assign _T_90 = _T_82[1:0]; // @[LZD.scala 44:32]
  assign _T_91 = _T_90 != 2'h0; // @[LZD.scala 39:14]
  assign _T_92 = _T_90[1]; // @[LZD.scala 39:21]
  assign _T_93 = _T_90[0]; // @[LZD.scala 39:30]
  assign _T_94 = ~ _T_93; // @[LZD.scala 39:27]
  assign _T_95 = _T_92 | _T_94; // @[LZD.scala 39:25]
  assign _T_96 = {_T_91,_T_95}; // @[Cat.scala 29:58]
  assign _T_97 = _T_89[1]; // @[Shift.scala 12:21]
  assign _T_98 = _T_96[1]; // @[Shift.scala 12:21]
  assign _T_99 = _T_97 | _T_98; // @[LZD.scala 49:16]
  assign _T_100 = ~ _T_98; // @[LZD.scala 49:27]
  assign _T_101 = _T_97 | _T_100; // @[LZD.scala 49:25]
  assign _T_102 = _T_89[0:0]; // @[LZD.scala 49:47]
  assign _T_103 = _T_96[0:0]; // @[LZD.scala 49:59]
  assign _T_104 = _T_97 ? _T_102 : _T_103; // @[LZD.scala 49:35]
  assign _T_106 = {_T_99,_T_101,_T_104}; // @[Cat.scala 29:58]
  assign _T_107 = _T_81[3:0]; // @[LZD.scala 44:32]
  assign _T_108 = _T_107[3:2]; // @[LZD.scala 43:32]
  assign _T_109 = _T_108 != 2'h0; // @[LZD.scala 39:14]
  assign _T_110 = _T_108[1]; // @[LZD.scala 39:21]
  assign _T_111 = _T_108[0]; // @[LZD.scala 39:30]
  assign _T_112 = ~ _T_111; // @[LZD.scala 39:27]
  assign _T_113 = _T_110 | _T_112; // @[LZD.scala 39:25]
  assign _T_114 = {_T_109,_T_113}; // @[Cat.scala 29:58]
  assign _T_115 = _T_107[1:0]; // @[LZD.scala 44:32]
  assign _T_116 = _T_115 != 2'h0; // @[LZD.scala 39:14]
  assign _T_117 = _T_115[1]; // @[LZD.scala 39:21]
  assign _T_118 = _T_115[0]; // @[LZD.scala 39:30]
  assign _T_119 = ~ _T_118; // @[LZD.scala 39:27]
  assign _T_120 = _T_117 | _T_119; // @[LZD.scala 39:25]
  assign _T_121 = {_T_116,_T_120}; // @[Cat.scala 29:58]
  assign _T_122 = _T_114[1]; // @[Shift.scala 12:21]
  assign _T_123 = _T_121[1]; // @[Shift.scala 12:21]
  assign _T_124 = _T_122 | _T_123; // @[LZD.scala 49:16]
  assign _T_125 = ~ _T_123; // @[LZD.scala 49:27]
  assign _T_126 = _T_122 | _T_125; // @[LZD.scala 49:25]
  assign _T_127 = _T_114[0:0]; // @[LZD.scala 49:47]
  assign _T_128 = _T_121[0:0]; // @[LZD.scala 49:59]
  assign _T_129 = _T_122 ? _T_127 : _T_128; // @[LZD.scala 49:35]
  assign _T_131 = {_T_124,_T_126,_T_129}; // @[Cat.scala 29:58]
  assign _T_132 = _T_106[2]; // @[Shift.scala 12:21]
  assign _T_133 = _T_131[2]; // @[Shift.scala 12:21]
  assign _T_134 = _T_132 | _T_133; // @[LZD.scala 49:16]
  assign _T_135 = ~ _T_133; // @[LZD.scala 49:27]
  assign _T_136 = _T_132 | _T_135; // @[LZD.scala 49:25]
  assign _T_137 = _T_106[1:0]; // @[LZD.scala 49:47]
  assign _T_138 = _T_131[1:0]; // @[LZD.scala 49:59]
  assign _T_139 = _T_132 ? _T_137 : _T_138; // @[LZD.scala 49:35]
  assign _T_141 = {_T_134,_T_136,_T_139}; // @[Cat.scala 29:58]
  assign _T_142 = _T_80[3]; // @[Shift.scala 12:21]
  assign _T_143 = _T_141[3]; // @[Shift.scala 12:21]
  assign _T_144 = _T_142 | _T_143; // @[LZD.scala 49:16]
  assign _T_145 = ~ _T_143; // @[LZD.scala 49:27]
  assign _T_146 = _T_142 | _T_145; // @[LZD.scala 49:25]
  assign _T_147 = _T_80[2:0]; // @[LZD.scala 49:47]
  assign _T_148 = _T_141[2:0]; // @[LZD.scala 49:59]
  assign _T_149 = _T_142 ? _T_147 : _T_148; // @[LZD.scala 49:35]
  assign _T_151 = {_T_144,_T_146,_T_149}; // @[Cat.scala 29:58]
  assign _T_152 = _T_18[12:0]; // @[LZD.scala 44:32]
  assign _T_153 = _T_152[12:5]; // @[LZD.scala 43:32]
  assign _T_154 = _T_153[7:4]; // @[LZD.scala 43:32]
  assign _T_155 = _T_154[3:2]; // @[LZD.scala 43:32]
  assign _T_156 = _T_155 != 2'h0; // @[LZD.scala 39:14]
  assign _T_157 = _T_155[1]; // @[LZD.scala 39:21]
  assign _T_158 = _T_155[0]; // @[LZD.scala 39:30]
  assign _T_159 = ~ _T_158; // @[LZD.scala 39:27]
  assign _T_160 = _T_157 | _T_159; // @[LZD.scala 39:25]
  assign _T_161 = {_T_156,_T_160}; // @[Cat.scala 29:58]
  assign _T_162 = _T_154[1:0]; // @[LZD.scala 44:32]
  assign _T_163 = _T_162 != 2'h0; // @[LZD.scala 39:14]
  assign _T_164 = _T_162[1]; // @[LZD.scala 39:21]
  assign _T_165 = _T_162[0]; // @[LZD.scala 39:30]
  assign _T_166 = ~ _T_165; // @[LZD.scala 39:27]
  assign _T_167 = _T_164 | _T_166; // @[LZD.scala 39:25]
  assign _T_168 = {_T_163,_T_167}; // @[Cat.scala 29:58]
  assign _T_169 = _T_161[1]; // @[Shift.scala 12:21]
  assign _T_170 = _T_168[1]; // @[Shift.scala 12:21]
  assign _T_171 = _T_169 | _T_170; // @[LZD.scala 49:16]
  assign _T_172 = ~ _T_170; // @[LZD.scala 49:27]
  assign _T_173 = _T_169 | _T_172; // @[LZD.scala 49:25]
  assign _T_174 = _T_161[0:0]; // @[LZD.scala 49:47]
  assign _T_175 = _T_168[0:0]; // @[LZD.scala 49:59]
  assign _T_176 = _T_169 ? _T_174 : _T_175; // @[LZD.scala 49:35]
  assign _T_178 = {_T_171,_T_173,_T_176}; // @[Cat.scala 29:58]
  assign _T_179 = _T_153[3:0]; // @[LZD.scala 44:32]
  assign _T_180 = _T_179[3:2]; // @[LZD.scala 43:32]
  assign _T_181 = _T_180 != 2'h0; // @[LZD.scala 39:14]
  assign _T_182 = _T_180[1]; // @[LZD.scala 39:21]
  assign _T_183 = _T_180[0]; // @[LZD.scala 39:30]
  assign _T_184 = ~ _T_183; // @[LZD.scala 39:27]
  assign _T_185 = _T_182 | _T_184; // @[LZD.scala 39:25]
  assign _T_186 = {_T_181,_T_185}; // @[Cat.scala 29:58]
  assign _T_187 = _T_179[1:0]; // @[LZD.scala 44:32]
  assign _T_188 = _T_187 != 2'h0; // @[LZD.scala 39:14]
  assign _T_189 = _T_187[1]; // @[LZD.scala 39:21]
  assign _T_190 = _T_187[0]; // @[LZD.scala 39:30]
  assign _T_191 = ~ _T_190; // @[LZD.scala 39:27]
  assign _T_192 = _T_189 | _T_191; // @[LZD.scala 39:25]
  assign _T_193 = {_T_188,_T_192}; // @[Cat.scala 29:58]
  assign _T_194 = _T_186[1]; // @[Shift.scala 12:21]
  assign _T_195 = _T_193[1]; // @[Shift.scala 12:21]
  assign _T_196 = _T_194 | _T_195; // @[LZD.scala 49:16]
  assign _T_197 = ~ _T_195; // @[LZD.scala 49:27]
  assign _T_198 = _T_194 | _T_197; // @[LZD.scala 49:25]
  assign _T_199 = _T_186[0:0]; // @[LZD.scala 49:47]
  assign _T_200 = _T_193[0:0]; // @[LZD.scala 49:59]
  assign _T_201 = _T_194 ? _T_199 : _T_200; // @[LZD.scala 49:35]
  assign _T_203 = {_T_196,_T_198,_T_201}; // @[Cat.scala 29:58]
  assign _T_204 = _T_178[2]; // @[Shift.scala 12:21]
  assign _T_205 = _T_203[2]; // @[Shift.scala 12:21]
  assign _T_206 = _T_204 | _T_205; // @[LZD.scala 49:16]
  assign _T_207 = ~ _T_205; // @[LZD.scala 49:27]
  assign _T_208 = _T_204 | _T_207; // @[LZD.scala 49:25]
  assign _T_209 = _T_178[1:0]; // @[LZD.scala 49:47]
  assign _T_210 = _T_203[1:0]; // @[LZD.scala 49:59]
  assign _T_211 = _T_204 ? _T_209 : _T_210; // @[LZD.scala 49:35]
  assign _T_213 = {_T_206,_T_208,_T_211}; // @[Cat.scala 29:58]
  assign _T_214 = _T_152[4:0]; // @[LZD.scala 44:32]
  assign _T_215 = _T_214[4:1]; // @[LZD.scala 43:32]
  assign _T_216 = _T_215[3:2]; // @[LZD.scala 43:32]
  assign _T_217 = _T_216 != 2'h0; // @[LZD.scala 39:14]
  assign _T_218 = _T_216[1]; // @[LZD.scala 39:21]
  assign _T_219 = _T_216[0]; // @[LZD.scala 39:30]
  assign _T_220 = ~ _T_219; // @[LZD.scala 39:27]
  assign _T_221 = _T_218 | _T_220; // @[LZD.scala 39:25]
  assign _T_222 = {_T_217,_T_221}; // @[Cat.scala 29:58]
  assign _T_223 = _T_215[1:0]; // @[LZD.scala 44:32]
  assign _T_224 = _T_223 != 2'h0; // @[LZD.scala 39:14]
  assign _T_225 = _T_223[1]; // @[LZD.scala 39:21]
  assign _T_226 = _T_223[0]; // @[LZD.scala 39:30]
  assign _T_227 = ~ _T_226; // @[LZD.scala 39:27]
  assign _T_228 = _T_225 | _T_227; // @[LZD.scala 39:25]
  assign _T_229 = {_T_224,_T_228}; // @[Cat.scala 29:58]
  assign _T_230 = _T_222[1]; // @[Shift.scala 12:21]
  assign _T_231 = _T_229[1]; // @[Shift.scala 12:21]
  assign _T_232 = _T_230 | _T_231; // @[LZD.scala 49:16]
  assign _T_233 = ~ _T_231; // @[LZD.scala 49:27]
  assign _T_234 = _T_230 | _T_233; // @[LZD.scala 49:25]
  assign _T_235 = _T_222[0:0]; // @[LZD.scala 49:47]
  assign _T_236 = _T_229[0:0]; // @[LZD.scala 49:59]
  assign _T_237 = _T_230 ? _T_235 : _T_236; // @[LZD.scala 49:35]
  assign _T_239 = {_T_232,_T_234,_T_237}; // @[Cat.scala 29:58]
  assign _T_240 = _T_214[0:0]; // @[LZD.scala 44:32]
  assign _T_242 = _T_239[2]; // @[Shift.scala 12:21]
  assign _T_244 = {1'h1,_T_240}; // @[Cat.scala 29:58]
  assign _T_245 = _T_239[1:0]; // @[LZD.scala 55:32]
  assign _T_246 = _T_242 ? _T_245 : _T_244; // @[LZD.scala 55:20]
  assign _T_247 = {_T_242,_T_246}; // @[Cat.scala 29:58]
  assign _T_248 = _T_213[3]; // @[Shift.scala 12:21]
  assign _T_250 = _T_213[2:0]; // @[LZD.scala 55:32]
  assign _T_251 = _T_248 ? _T_250 : _T_247; // @[LZD.scala 55:20]
  assign _T_252 = {_T_248,_T_251}; // @[Cat.scala 29:58]
  assign _T_253 = _T_151[4]; // @[Shift.scala 12:21]
  assign _T_255 = _T_151[3:0]; // @[LZD.scala 55:32]
  assign _T_256 = _T_253 ? _T_255 : _T_252; // @[LZD.scala 55:20]
  assign _T_257 = {_T_253,_T_256}; // @[Cat.scala 29:58]
  assign _T_258 = ~ _T_257; // @[convert.scala 21:22]
  assign _T_259 = realA[27:0]; // @[convert.scala 22:36]
  assign _T_260 = _T_258 < 5'h1c; // @[Shift.scala 16:24]
  assign _T_262 = _T_258[4]; // @[Shift.scala 12:21]
  assign _T_263 = _T_259[11:0]; // @[Shift.scala 64:52]
  assign _T_265 = {_T_263,16'h0}; // @[Cat.scala 29:58]
  assign _T_266 = _T_262 ? _T_265 : _T_259; // @[Shift.scala 64:27]
  assign _T_267 = _T_258[3:0]; // @[Shift.scala 66:70]
  assign _T_268 = _T_267[3]; // @[Shift.scala 12:21]
  assign _T_269 = _T_266[19:0]; // @[Shift.scala 64:52]
  assign _T_271 = {_T_269,8'h0}; // @[Cat.scala 29:58]
  assign _T_272 = _T_268 ? _T_271 : _T_266; // @[Shift.scala 64:27]
  assign _T_273 = _T_267[2:0]; // @[Shift.scala 66:70]
  assign _T_274 = _T_273[2]; // @[Shift.scala 12:21]
  assign _T_275 = _T_272[23:0]; // @[Shift.scala 64:52]
  assign _T_277 = {_T_275,4'h0}; // @[Cat.scala 29:58]
  assign _T_278 = _T_274 ? _T_277 : _T_272; // @[Shift.scala 64:27]
  assign _T_279 = _T_273[1:0]; // @[Shift.scala 66:70]
  assign _T_280 = _T_279[1]; // @[Shift.scala 12:21]
  assign _T_281 = _T_278[25:0]; // @[Shift.scala 64:52]
  assign _T_283 = {_T_281,2'h0}; // @[Cat.scala 29:58]
  assign _T_284 = _T_280 ? _T_283 : _T_278; // @[Shift.scala 64:27]
  assign _T_285 = _T_279[0:0]; // @[Shift.scala 66:70]
  assign _T_287 = _T_284[26:0]; // @[Shift.scala 64:52]
  assign _T_288 = {_T_287,1'h0}; // @[Cat.scala 29:58]
  assign _T_289 = _T_285 ? _T_288 : _T_284; // @[Shift.scala 64:27]
  assign _T_290 = _T_260 ? _T_289 : 28'h0; // @[Shift.scala 16:10]
  assign _T_291 = _T_290[27:25]; // @[convert.scala 23:34]
  assign decA_fraction = _T_290[24:0]; // @[convert.scala 24:34]
  assign _T_293 = _T_15 == 1'h0; // @[convert.scala 25:26]
  assign _T_295 = _T_15 ? _T_258 : _T_257; // @[convert.scala 25:42]
  assign _T_298 = ~ _T_291; // @[convert.scala 26:67]
  assign _T_299 = _T_13 ? _T_298 : _T_291; // @[convert.scala 26:51]
  assign _T_300 = {_T_293,_T_295,_T_299}; // @[Cat.scala 29:58]
  assign _T_302 = realA[29:0]; // @[convert.scala 29:56]
  assign _T_303 = _T_302 != 30'h0; // @[convert.scala 29:60]
  assign _T_304 = ~ _T_303; // @[convert.scala 29:41]
  assign decA_isNaR = _T_13 & _T_304; // @[convert.scala 29:39]
  assign _T_307 = _T_13 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_307 & _T_304; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_300); // @[convert.scala 32:24]
  assign _T_316 = io_B[30]; // @[convert.scala 18:24]
  assign _T_317 = io_B[29]; // @[convert.scala 18:40]
  assign _T_318 = _T_316 ^ _T_317; // @[convert.scala 18:36]
  assign _T_319 = io_B[29:1]; // @[convert.scala 19:24]
  assign _T_320 = io_B[28:0]; // @[convert.scala 19:43]
  assign _T_321 = _T_319 ^ _T_320; // @[convert.scala 19:39]
  assign _T_322 = _T_321[28:13]; // @[LZD.scala 43:32]
  assign _T_323 = _T_322[15:8]; // @[LZD.scala 43:32]
  assign _T_324 = _T_323[7:4]; // @[LZD.scala 43:32]
  assign _T_325 = _T_324[3:2]; // @[LZD.scala 43:32]
  assign _T_326 = _T_325 != 2'h0; // @[LZD.scala 39:14]
  assign _T_327 = _T_325[1]; // @[LZD.scala 39:21]
  assign _T_328 = _T_325[0]; // @[LZD.scala 39:30]
  assign _T_329 = ~ _T_328; // @[LZD.scala 39:27]
  assign _T_330 = _T_327 | _T_329; // @[LZD.scala 39:25]
  assign _T_331 = {_T_326,_T_330}; // @[Cat.scala 29:58]
  assign _T_332 = _T_324[1:0]; // @[LZD.scala 44:32]
  assign _T_333 = _T_332 != 2'h0; // @[LZD.scala 39:14]
  assign _T_334 = _T_332[1]; // @[LZD.scala 39:21]
  assign _T_335 = _T_332[0]; // @[LZD.scala 39:30]
  assign _T_336 = ~ _T_335; // @[LZD.scala 39:27]
  assign _T_337 = _T_334 | _T_336; // @[LZD.scala 39:25]
  assign _T_338 = {_T_333,_T_337}; // @[Cat.scala 29:58]
  assign _T_339 = _T_331[1]; // @[Shift.scala 12:21]
  assign _T_340 = _T_338[1]; // @[Shift.scala 12:21]
  assign _T_341 = _T_339 | _T_340; // @[LZD.scala 49:16]
  assign _T_342 = ~ _T_340; // @[LZD.scala 49:27]
  assign _T_343 = _T_339 | _T_342; // @[LZD.scala 49:25]
  assign _T_344 = _T_331[0:0]; // @[LZD.scala 49:47]
  assign _T_345 = _T_338[0:0]; // @[LZD.scala 49:59]
  assign _T_346 = _T_339 ? _T_344 : _T_345; // @[LZD.scala 49:35]
  assign _T_348 = {_T_341,_T_343,_T_346}; // @[Cat.scala 29:58]
  assign _T_349 = _T_323[3:0]; // @[LZD.scala 44:32]
  assign _T_350 = _T_349[3:2]; // @[LZD.scala 43:32]
  assign _T_351 = _T_350 != 2'h0; // @[LZD.scala 39:14]
  assign _T_352 = _T_350[1]; // @[LZD.scala 39:21]
  assign _T_353 = _T_350[0]; // @[LZD.scala 39:30]
  assign _T_354 = ~ _T_353; // @[LZD.scala 39:27]
  assign _T_355 = _T_352 | _T_354; // @[LZD.scala 39:25]
  assign _T_356 = {_T_351,_T_355}; // @[Cat.scala 29:58]
  assign _T_357 = _T_349[1:0]; // @[LZD.scala 44:32]
  assign _T_358 = _T_357 != 2'h0; // @[LZD.scala 39:14]
  assign _T_359 = _T_357[1]; // @[LZD.scala 39:21]
  assign _T_360 = _T_357[0]; // @[LZD.scala 39:30]
  assign _T_361 = ~ _T_360; // @[LZD.scala 39:27]
  assign _T_362 = _T_359 | _T_361; // @[LZD.scala 39:25]
  assign _T_363 = {_T_358,_T_362}; // @[Cat.scala 29:58]
  assign _T_364 = _T_356[1]; // @[Shift.scala 12:21]
  assign _T_365 = _T_363[1]; // @[Shift.scala 12:21]
  assign _T_366 = _T_364 | _T_365; // @[LZD.scala 49:16]
  assign _T_367 = ~ _T_365; // @[LZD.scala 49:27]
  assign _T_368 = _T_364 | _T_367; // @[LZD.scala 49:25]
  assign _T_369 = _T_356[0:0]; // @[LZD.scala 49:47]
  assign _T_370 = _T_363[0:0]; // @[LZD.scala 49:59]
  assign _T_371 = _T_364 ? _T_369 : _T_370; // @[LZD.scala 49:35]
  assign _T_373 = {_T_366,_T_368,_T_371}; // @[Cat.scala 29:58]
  assign _T_374 = _T_348[2]; // @[Shift.scala 12:21]
  assign _T_375 = _T_373[2]; // @[Shift.scala 12:21]
  assign _T_376 = _T_374 | _T_375; // @[LZD.scala 49:16]
  assign _T_377 = ~ _T_375; // @[LZD.scala 49:27]
  assign _T_378 = _T_374 | _T_377; // @[LZD.scala 49:25]
  assign _T_379 = _T_348[1:0]; // @[LZD.scala 49:47]
  assign _T_380 = _T_373[1:0]; // @[LZD.scala 49:59]
  assign _T_381 = _T_374 ? _T_379 : _T_380; // @[LZD.scala 49:35]
  assign _T_383 = {_T_376,_T_378,_T_381}; // @[Cat.scala 29:58]
  assign _T_384 = _T_322[7:0]; // @[LZD.scala 44:32]
  assign _T_385 = _T_384[7:4]; // @[LZD.scala 43:32]
  assign _T_386 = _T_385[3:2]; // @[LZD.scala 43:32]
  assign _T_387 = _T_386 != 2'h0; // @[LZD.scala 39:14]
  assign _T_388 = _T_386[1]; // @[LZD.scala 39:21]
  assign _T_389 = _T_386[0]; // @[LZD.scala 39:30]
  assign _T_390 = ~ _T_389; // @[LZD.scala 39:27]
  assign _T_391 = _T_388 | _T_390; // @[LZD.scala 39:25]
  assign _T_392 = {_T_387,_T_391}; // @[Cat.scala 29:58]
  assign _T_393 = _T_385[1:0]; // @[LZD.scala 44:32]
  assign _T_394 = _T_393 != 2'h0; // @[LZD.scala 39:14]
  assign _T_395 = _T_393[1]; // @[LZD.scala 39:21]
  assign _T_396 = _T_393[0]; // @[LZD.scala 39:30]
  assign _T_397 = ~ _T_396; // @[LZD.scala 39:27]
  assign _T_398 = _T_395 | _T_397; // @[LZD.scala 39:25]
  assign _T_399 = {_T_394,_T_398}; // @[Cat.scala 29:58]
  assign _T_400 = _T_392[1]; // @[Shift.scala 12:21]
  assign _T_401 = _T_399[1]; // @[Shift.scala 12:21]
  assign _T_402 = _T_400 | _T_401; // @[LZD.scala 49:16]
  assign _T_403 = ~ _T_401; // @[LZD.scala 49:27]
  assign _T_404 = _T_400 | _T_403; // @[LZD.scala 49:25]
  assign _T_405 = _T_392[0:0]; // @[LZD.scala 49:47]
  assign _T_406 = _T_399[0:0]; // @[LZD.scala 49:59]
  assign _T_407 = _T_400 ? _T_405 : _T_406; // @[LZD.scala 49:35]
  assign _T_409 = {_T_402,_T_404,_T_407}; // @[Cat.scala 29:58]
  assign _T_410 = _T_384[3:0]; // @[LZD.scala 44:32]
  assign _T_411 = _T_410[3:2]; // @[LZD.scala 43:32]
  assign _T_412 = _T_411 != 2'h0; // @[LZD.scala 39:14]
  assign _T_413 = _T_411[1]; // @[LZD.scala 39:21]
  assign _T_414 = _T_411[0]; // @[LZD.scala 39:30]
  assign _T_415 = ~ _T_414; // @[LZD.scala 39:27]
  assign _T_416 = _T_413 | _T_415; // @[LZD.scala 39:25]
  assign _T_417 = {_T_412,_T_416}; // @[Cat.scala 29:58]
  assign _T_418 = _T_410[1:0]; // @[LZD.scala 44:32]
  assign _T_419 = _T_418 != 2'h0; // @[LZD.scala 39:14]
  assign _T_420 = _T_418[1]; // @[LZD.scala 39:21]
  assign _T_421 = _T_418[0]; // @[LZD.scala 39:30]
  assign _T_422 = ~ _T_421; // @[LZD.scala 39:27]
  assign _T_423 = _T_420 | _T_422; // @[LZD.scala 39:25]
  assign _T_424 = {_T_419,_T_423}; // @[Cat.scala 29:58]
  assign _T_425 = _T_417[1]; // @[Shift.scala 12:21]
  assign _T_426 = _T_424[1]; // @[Shift.scala 12:21]
  assign _T_427 = _T_425 | _T_426; // @[LZD.scala 49:16]
  assign _T_428 = ~ _T_426; // @[LZD.scala 49:27]
  assign _T_429 = _T_425 | _T_428; // @[LZD.scala 49:25]
  assign _T_430 = _T_417[0:0]; // @[LZD.scala 49:47]
  assign _T_431 = _T_424[0:0]; // @[LZD.scala 49:59]
  assign _T_432 = _T_425 ? _T_430 : _T_431; // @[LZD.scala 49:35]
  assign _T_434 = {_T_427,_T_429,_T_432}; // @[Cat.scala 29:58]
  assign _T_435 = _T_409[2]; // @[Shift.scala 12:21]
  assign _T_436 = _T_434[2]; // @[Shift.scala 12:21]
  assign _T_437 = _T_435 | _T_436; // @[LZD.scala 49:16]
  assign _T_438 = ~ _T_436; // @[LZD.scala 49:27]
  assign _T_439 = _T_435 | _T_438; // @[LZD.scala 49:25]
  assign _T_440 = _T_409[1:0]; // @[LZD.scala 49:47]
  assign _T_441 = _T_434[1:0]; // @[LZD.scala 49:59]
  assign _T_442 = _T_435 ? _T_440 : _T_441; // @[LZD.scala 49:35]
  assign _T_444 = {_T_437,_T_439,_T_442}; // @[Cat.scala 29:58]
  assign _T_445 = _T_383[3]; // @[Shift.scala 12:21]
  assign _T_446 = _T_444[3]; // @[Shift.scala 12:21]
  assign _T_447 = _T_445 | _T_446; // @[LZD.scala 49:16]
  assign _T_448 = ~ _T_446; // @[LZD.scala 49:27]
  assign _T_449 = _T_445 | _T_448; // @[LZD.scala 49:25]
  assign _T_450 = _T_383[2:0]; // @[LZD.scala 49:47]
  assign _T_451 = _T_444[2:0]; // @[LZD.scala 49:59]
  assign _T_452 = _T_445 ? _T_450 : _T_451; // @[LZD.scala 49:35]
  assign _T_454 = {_T_447,_T_449,_T_452}; // @[Cat.scala 29:58]
  assign _T_455 = _T_321[12:0]; // @[LZD.scala 44:32]
  assign _T_456 = _T_455[12:5]; // @[LZD.scala 43:32]
  assign _T_457 = _T_456[7:4]; // @[LZD.scala 43:32]
  assign _T_458 = _T_457[3:2]; // @[LZD.scala 43:32]
  assign _T_459 = _T_458 != 2'h0; // @[LZD.scala 39:14]
  assign _T_460 = _T_458[1]; // @[LZD.scala 39:21]
  assign _T_461 = _T_458[0]; // @[LZD.scala 39:30]
  assign _T_462 = ~ _T_461; // @[LZD.scala 39:27]
  assign _T_463 = _T_460 | _T_462; // @[LZD.scala 39:25]
  assign _T_464 = {_T_459,_T_463}; // @[Cat.scala 29:58]
  assign _T_465 = _T_457[1:0]; // @[LZD.scala 44:32]
  assign _T_466 = _T_465 != 2'h0; // @[LZD.scala 39:14]
  assign _T_467 = _T_465[1]; // @[LZD.scala 39:21]
  assign _T_468 = _T_465[0]; // @[LZD.scala 39:30]
  assign _T_469 = ~ _T_468; // @[LZD.scala 39:27]
  assign _T_470 = _T_467 | _T_469; // @[LZD.scala 39:25]
  assign _T_471 = {_T_466,_T_470}; // @[Cat.scala 29:58]
  assign _T_472 = _T_464[1]; // @[Shift.scala 12:21]
  assign _T_473 = _T_471[1]; // @[Shift.scala 12:21]
  assign _T_474 = _T_472 | _T_473; // @[LZD.scala 49:16]
  assign _T_475 = ~ _T_473; // @[LZD.scala 49:27]
  assign _T_476 = _T_472 | _T_475; // @[LZD.scala 49:25]
  assign _T_477 = _T_464[0:0]; // @[LZD.scala 49:47]
  assign _T_478 = _T_471[0:0]; // @[LZD.scala 49:59]
  assign _T_479 = _T_472 ? _T_477 : _T_478; // @[LZD.scala 49:35]
  assign _T_481 = {_T_474,_T_476,_T_479}; // @[Cat.scala 29:58]
  assign _T_482 = _T_456[3:0]; // @[LZD.scala 44:32]
  assign _T_483 = _T_482[3:2]; // @[LZD.scala 43:32]
  assign _T_484 = _T_483 != 2'h0; // @[LZD.scala 39:14]
  assign _T_485 = _T_483[1]; // @[LZD.scala 39:21]
  assign _T_486 = _T_483[0]; // @[LZD.scala 39:30]
  assign _T_487 = ~ _T_486; // @[LZD.scala 39:27]
  assign _T_488 = _T_485 | _T_487; // @[LZD.scala 39:25]
  assign _T_489 = {_T_484,_T_488}; // @[Cat.scala 29:58]
  assign _T_490 = _T_482[1:0]; // @[LZD.scala 44:32]
  assign _T_491 = _T_490 != 2'h0; // @[LZD.scala 39:14]
  assign _T_492 = _T_490[1]; // @[LZD.scala 39:21]
  assign _T_493 = _T_490[0]; // @[LZD.scala 39:30]
  assign _T_494 = ~ _T_493; // @[LZD.scala 39:27]
  assign _T_495 = _T_492 | _T_494; // @[LZD.scala 39:25]
  assign _T_496 = {_T_491,_T_495}; // @[Cat.scala 29:58]
  assign _T_497 = _T_489[1]; // @[Shift.scala 12:21]
  assign _T_498 = _T_496[1]; // @[Shift.scala 12:21]
  assign _T_499 = _T_497 | _T_498; // @[LZD.scala 49:16]
  assign _T_500 = ~ _T_498; // @[LZD.scala 49:27]
  assign _T_501 = _T_497 | _T_500; // @[LZD.scala 49:25]
  assign _T_502 = _T_489[0:0]; // @[LZD.scala 49:47]
  assign _T_503 = _T_496[0:0]; // @[LZD.scala 49:59]
  assign _T_504 = _T_497 ? _T_502 : _T_503; // @[LZD.scala 49:35]
  assign _T_506 = {_T_499,_T_501,_T_504}; // @[Cat.scala 29:58]
  assign _T_507 = _T_481[2]; // @[Shift.scala 12:21]
  assign _T_508 = _T_506[2]; // @[Shift.scala 12:21]
  assign _T_509 = _T_507 | _T_508; // @[LZD.scala 49:16]
  assign _T_510 = ~ _T_508; // @[LZD.scala 49:27]
  assign _T_511 = _T_507 | _T_510; // @[LZD.scala 49:25]
  assign _T_512 = _T_481[1:0]; // @[LZD.scala 49:47]
  assign _T_513 = _T_506[1:0]; // @[LZD.scala 49:59]
  assign _T_514 = _T_507 ? _T_512 : _T_513; // @[LZD.scala 49:35]
  assign _T_516 = {_T_509,_T_511,_T_514}; // @[Cat.scala 29:58]
  assign _T_517 = _T_455[4:0]; // @[LZD.scala 44:32]
  assign _T_518 = _T_517[4:1]; // @[LZD.scala 43:32]
  assign _T_519 = _T_518[3:2]; // @[LZD.scala 43:32]
  assign _T_520 = _T_519 != 2'h0; // @[LZD.scala 39:14]
  assign _T_521 = _T_519[1]; // @[LZD.scala 39:21]
  assign _T_522 = _T_519[0]; // @[LZD.scala 39:30]
  assign _T_523 = ~ _T_522; // @[LZD.scala 39:27]
  assign _T_524 = _T_521 | _T_523; // @[LZD.scala 39:25]
  assign _T_525 = {_T_520,_T_524}; // @[Cat.scala 29:58]
  assign _T_526 = _T_518[1:0]; // @[LZD.scala 44:32]
  assign _T_527 = _T_526 != 2'h0; // @[LZD.scala 39:14]
  assign _T_528 = _T_526[1]; // @[LZD.scala 39:21]
  assign _T_529 = _T_526[0]; // @[LZD.scala 39:30]
  assign _T_530 = ~ _T_529; // @[LZD.scala 39:27]
  assign _T_531 = _T_528 | _T_530; // @[LZD.scala 39:25]
  assign _T_532 = {_T_527,_T_531}; // @[Cat.scala 29:58]
  assign _T_533 = _T_525[1]; // @[Shift.scala 12:21]
  assign _T_534 = _T_532[1]; // @[Shift.scala 12:21]
  assign _T_535 = _T_533 | _T_534; // @[LZD.scala 49:16]
  assign _T_536 = ~ _T_534; // @[LZD.scala 49:27]
  assign _T_537 = _T_533 | _T_536; // @[LZD.scala 49:25]
  assign _T_538 = _T_525[0:0]; // @[LZD.scala 49:47]
  assign _T_539 = _T_532[0:0]; // @[LZD.scala 49:59]
  assign _T_540 = _T_533 ? _T_538 : _T_539; // @[LZD.scala 49:35]
  assign _T_542 = {_T_535,_T_537,_T_540}; // @[Cat.scala 29:58]
  assign _T_543 = _T_517[0:0]; // @[LZD.scala 44:32]
  assign _T_545 = _T_542[2]; // @[Shift.scala 12:21]
  assign _T_547 = {1'h1,_T_543}; // @[Cat.scala 29:58]
  assign _T_548 = _T_542[1:0]; // @[LZD.scala 55:32]
  assign _T_549 = _T_545 ? _T_548 : _T_547; // @[LZD.scala 55:20]
  assign _T_550 = {_T_545,_T_549}; // @[Cat.scala 29:58]
  assign _T_551 = _T_516[3]; // @[Shift.scala 12:21]
  assign _T_553 = _T_516[2:0]; // @[LZD.scala 55:32]
  assign _T_554 = _T_551 ? _T_553 : _T_550; // @[LZD.scala 55:20]
  assign _T_555 = {_T_551,_T_554}; // @[Cat.scala 29:58]
  assign _T_556 = _T_454[4]; // @[Shift.scala 12:21]
  assign _T_558 = _T_454[3:0]; // @[LZD.scala 55:32]
  assign _T_559 = _T_556 ? _T_558 : _T_555; // @[LZD.scala 55:20]
  assign _T_560 = {_T_556,_T_559}; // @[Cat.scala 29:58]
  assign _T_561 = ~ _T_560; // @[convert.scala 21:22]
  assign _T_562 = io_B[27:0]; // @[convert.scala 22:36]
  assign _T_563 = _T_561 < 5'h1c; // @[Shift.scala 16:24]
  assign _T_565 = _T_561[4]; // @[Shift.scala 12:21]
  assign _T_566 = _T_562[11:0]; // @[Shift.scala 64:52]
  assign _T_568 = {_T_566,16'h0}; // @[Cat.scala 29:58]
  assign _T_569 = _T_565 ? _T_568 : _T_562; // @[Shift.scala 64:27]
  assign _T_570 = _T_561[3:0]; // @[Shift.scala 66:70]
  assign _T_571 = _T_570[3]; // @[Shift.scala 12:21]
  assign _T_572 = _T_569[19:0]; // @[Shift.scala 64:52]
  assign _T_574 = {_T_572,8'h0}; // @[Cat.scala 29:58]
  assign _T_575 = _T_571 ? _T_574 : _T_569; // @[Shift.scala 64:27]
  assign _T_576 = _T_570[2:0]; // @[Shift.scala 66:70]
  assign _T_577 = _T_576[2]; // @[Shift.scala 12:21]
  assign _T_578 = _T_575[23:0]; // @[Shift.scala 64:52]
  assign _T_580 = {_T_578,4'h0}; // @[Cat.scala 29:58]
  assign _T_581 = _T_577 ? _T_580 : _T_575; // @[Shift.scala 64:27]
  assign _T_582 = _T_576[1:0]; // @[Shift.scala 66:70]
  assign _T_583 = _T_582[1]; // @[Shift.scala 12:21]
  assign _T_584 = _T_581[25:0]; // @[Shift.scala 64:52]
  assign _T_586 = {_T_584,2'h0}; // @[Cat.scala 29:58]
  assign _T_587 = _T_583 ? _T_586 : _T_581; // @[Shift.scala 64:27]
  assign _T_588 = _T_582[0:0]; // @[Shift.scala 66:70]
  assign _T_590 = _T_587[26:0]; // @[Shift.scala 64:52]
  assign _T_591 = {_T_590,1'h0}; // @[Cat.scala 29:58]
  assign _T_592 = _T_588 ? _T_591 : _T_587; // @[Shift.scala 64:27]
  assign _T_593 = _T_563 ? _T_592 : 28'h0; // @[Shift.scala 16:10]
  assign _T_594 = _T_593[27:25]; // @[convert.scala 23:34]
  assign decB_fraction = _T_593[24:0]; // @[convert.scala 24:34]
  assign _T_596 = _T_318 == 1'h0; // @[convert.scala 25:26]
  assign _T_598 = _T_318 ? _T_561 : _T_560; // @[convert.scala 25:42]
  assign _T_601 = ~ _T_594; // @[convert.scala 26:67]
  assign _T_602 = _T_316 ? _T_601 : _T_594; // @[convert.scala 26:51]
  assign _T_603 = {_T_596,_T_598,_T_602}; // @[Cat.scala 29:58]
  assign _T_605 = io_B[29:0]; // @[convert.scala 29:56]
  assign _T_606 = _T_605 != 30'h0; // @[convert.scala 29:60]
  assign _T_607 = ~ _T_606; // @[convert.scala 29:41]
  assign decB_isNaR = _T_316 & _T_607; // @[convert.scala 29:39]
  assign _T_610 = _T_316 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_610 & _T_607; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_603); // @[convert.scala 32:24]
  assign _T_619 = realC[30]; // @[convert.scala 18:24]
  assign _T_620 = realC[29]; // @[convert.scala 18:40]
  assign _T_621 = _T_619 ^ _T_620; // @[convert.scala 18:36]
  assign _T_622 = realC[29:1]; // @[convert.scala 19:24]
  assign _T_623 = realC[28:0]; // @[convert.scala 19:43]
  assign _T_624 = _T_622 ^ _T_623; // @[convert.scala 19:39]
  assign _T_625 = _T_624[28:13]; // @[LZD.scala 43:32]
  assign _T_626 = _T_625[15:8]; // @[LZD.scala 43:32]
  assign _T_627 = _T_626[7:4]; // @[LZD.scala 43:32]
  assign _T_628 = _T_627[3:2]; // @[LZD.scala 43:32]
  assign _T_629 = _T_628 != 2'h0; // @[LZD.scala 39:14]
  assign _T_630 = _T_628[1]; // @[LZD.scala 39:21]
  assign _T_631 = _T_628[0]; // @[LZD.scala 39:30]
  assign _T_632 = ~ _T_631; // @[LZD.scala 39:27]
  assign _T_633 = _T_630 | _T_632; // @[LZD.scala 39:25]
  assign _T_634 = {_T_629,_T_633}; // @[Cat.scala 29:58]
  assign _T_635 = _T_627[1:0]; // @[LZD.scala 44:32]
  assign _T_636 = _T_635 != 2'h0; // @[LZD.scala 39:14]
  assign _T_637 = _T_635[1]; // @[LZD.scala 39:21]
  assign _T_638 = _T_635[0]; // @[LZD.scala 39:30]
  assign _T_639 = ~ _T_638; // @[LZD.scala 39:27]
  assign _T_640 = _T_637 | _T_639; // @[LZD.scala 39:25]
  assign _T_641 = {_T_636,_T_640}; // @[Cat.scala 29:58]
  assign _T_642 = _T_634[1]; // @[Shift.scala 12:21]
  assign _T_643 = _T_641[1]; // @[Shift.scala 12:21]
  assign _T_644 = _T_642 | _T_643; // @[LZD.scala 49:16]
  assign _T_645 = ~ _T_643; // @[LZD.scala 49:27]
  assign _T_646 = _T_642 | _T_645; // @[LZD.scala 49:25]
  assign _T_647 = _T_634[0:0]; // @[LZD.scala 49:47]
  assign _T_648 = _T_641[0:0]; // @[LZD.scala 49:59]
  assign _T_649 = _T_642 ? _T_647 : _T_648; // @[LZD.scala 49:35]
  assign _T_651 = {_T_644,_T_646,_T_649}; // @[Cat.scala 29:58]
  assign _T_652 = _T_626[3:0]; // @[LZD.scala 44:32]
  assign _T_653 = _T_652[3:2]; // @[LZD.scala 43:32]
  assign _T_654 = _T_653 != 2'h0; // @[LZD.scala 39:14]
  assign _T_655 = _T_653[1]; // @[LZD.scala 39:21]
  assign _T_656 = _T_653[0]; // @[LZD.scala 39:30]
  assign _T_657 = ~ _T_656; // @[LZD.scala 39:27]
  assign _T_658 = _T_655 | _T_657; // @[LZD.scala 39:25]
  assign _T_659 = {_T_654,_T_658}; // @[Cat.scala 29:58]
  assign _T_660 = _T_652[1:0]; // @[LZD.scala 44:32]
  assign _T_661 = _T_660 != 2'h0; // @[LZD.scala 39:14]
  assign _T_662 = _T_660[1]; // @[LZD.scala 39:21]
  assign _T_663 = _T_660[0]; // @[LZD.scala 39:30]
  assign _T_664 = ~ _T_663; // @[LZD.scala 39:27]
  assign _T_665 = _T_662 | _T_664; // @[LZD.scala 39:25]
  assign _T_666 = {_T_661,_T_665}; // @[Cat.scala 29:58]
  assign _T_667 = _T_659[1]; // @[Shift.scala 12:21]
  assign _T_668 = _T_666[1]; // @[Shift.scala 12:21]
  assign _T_669 = _T_667 | _T_668; // @[LZD.scala 49:16]
  assign _T_670 = ~ _T_668; // @[LZD.scala 49:27]
  assign _T_671 = _T_667 | _T_670; // @[LZD.scala 49:25]
  assign _T_672 = _T_659[0:0]; // @[LZD.scala 49:47]
  assign _T_673 = _T_666[0:0]; // @[LZD.scala 49:59]
  assign _T_674 = _T_667 ? _T_672 : _T_673; // @[LZD.scala 49:35]
  assign _T_676 = {_T_669,_T_671,_T_674}; // @[Cat.scala 29:58]
  assign _T_677 = _T_651[2]; // @[Shift.scala 12:21]
  assign _T_678 = _T_676[2]; // @[Shift.scala 12:21]
  assign _T_679 = _T_677 | _T_678; // @[LZD.scala 49:16]
  assign _T_680 = ~ _T_678; // @[LZD.scala 49:27]
  assign _T_681 = _T_677 | _T_680; // @[LZD.scala 49:25]
  assign _T_682 = _T_651[1:0]; // @[LZD.scala 49:47]
  assign _T_683 = _T_676[1:0]; // @[LZD.scala 49:59]
  assign _T_684 = _T_677 ? _T_682 : _T_683; // @[LZD.scala 49:35]
  assign _T_686 = {_T_679,_T_681,_T_684}; // @[Cat.scala 29:58]
  assign _T_687 = _T_625[7:0]; // @[LZD.scala 44:32]
  assign _T_688 = _T_687[7:4]; // @[LZD.scala 43:32]
  assign _T_689 = _T_688[3:2]; // @[LZD.scala 43:32]
  assign _T_690 = _T_689 != 2'h0; // @[LZD.scala 39:14]
  assign _T_691 = _T_689[1]; // @[LZD.scala 39:21]
  assign _T_692 = _T_689[0]; // @[LZD.scala 39:30]
  assign _T_693 = ~ _T_692; // @[LZD.scala 39:27]
  assign _T_694 = _T_691 | _T_693; // @[LZD.scala 39:25]
  assign _T_695 = {_T_690,_T_694}; // @[Cat.scala 29:58]
  assign _T_696 = _T_688[1:0]; // @[LZD.scala 44:32]
  assign _T_697 = _T_696 != 2'h0; // @[LZD.scala 39:14]
  assign _T_698 = _T_696[1]; // @[LZD.scala 39:21]
  assign _T_699 = _T_696[0]; // @[LZD.scala 39:30]
  assign _T_700 = ~ _T_699; // @[LZD.scala 39:27]
  assign _T_701 = _T_698 | _T_700; // @[LZD.scala 39:25]
  assign _T_702 = {_T_697,_T_701}; // @[Cat.scala 29:58]
  assign _T_703 = _T_695[1]; // @[Shift.scala 12:21]
  assign _T_704 = _T_702[1]; // @[Shift.scala 12:21]
  assign _T_705 = _T_703 | _T_704; // @[LZD.scala 49:16]
  assign _T_706 = ~ _T_704; // @[LZD.scala 49:27]
  assign _T_707 = _T_703 | _T_706; // @[LZD.scala 49:25]
  assign _T_708 = _T_695[0:0]; // @[LZD.scala 49:47]
  assign _T_709 = _T_702[0:0]; // @[LZD.scala 49:59]
  assign _T_710 = _T_703 ? _T_708 : _T_709; // @[LZD.scala 49:35]
  assign _T_712 = {_T_705,_T_707,_T_710}; // @[Cat.scala 29:58]
  assign _T_713 = _T_687[3:0]; // @[LZD.scala 44:32]
  assign _T_714 = _T_713[3:2]; // @[LZD.scala 43:32]
  assign _T_715 = _T_714 != 2'h0; // @[LZD.scala 39:14]
  assign _T_716 = _T_714[1]; // @[LZD.scala 39:21]
  assign _T_717 = _T_714[0]; // @[LZD.scala 39:30]
  assign _T_718 = ~ _T_717; // @[LZD.scala 39:27]
  assign _T_719 = _T_716 | _T_718; // @[LZD.scala 39:25]
  assign _T_720 = {_T_715,_T_719}; // @[Cat.scala 29:58]
  assign _T_721 = _T_713[1:0]; // @[LZD.scala 44:32]
  assign _T_722 = _T_721 != 2'h0; // @[LZD.scala 39:14]
  assign _T_723 = _T_721[1]; // @[LZD.scala 39:21]
  assign _T_724 = _T_721[0]; // @[LZD.scala 39:30]
  assign _T_725 = ~ _T_724; // @[LZD.scala 39:27]
  assign _T_726 = _T_723 | _T_725; // @[LZD.scala 39:25]
  assign _T_727 = {_T_722,_T_726}; // @[Cat.scala 29:58]
  assign _T_728 = _T_720[1]; // @[Shift.scala 12:21]
  assign _T_729 = _T_727[1]; // @[Shift.scala 12:21]
  assign _T_730 = _T_728 | _T_729; // @[LZD.scala 49:16]
  assign _T_731 = ~ _T_729; // @[LZD.scala 49:27]
  assign _T_732 = _T_728 | _T_731; // @[LZD.scala 49:25]
  assign _T_733 = _T_720[0:0]; // @[LZD.scala 49:47]
  assign _T_734 = _T_727[0:0]; // @[LZD.scala 49:59]
  assign _T_735 = _T_728 ? _T_733 : _T_734; // @[LZD.scala 49:35]
  assign _T_737 = {_T_730,_T_732,_T_735}; // @[Cat.scala 29:58]
  assign _T_738 = _T_712[2]; // @[Shift.scala 12:21]
  assign _T_739 = _T_737[2]; // @[Shift.scala 12:21]
  assign _T_740 = _T_738 | _T_739; // @[LZD.scala 49:16]
  assign _T_741 = ~ _T_739; // @[LZD.scala 49:27]
  assign _T_742 = _T_738 | _T_741; // @[LZD.scala 49:25]
  assign _T_743 = _T_712[1:0]; // @[LZD.scala 49:47]
  assign _T_744 = _T_737[1:0]; // @[LZD.scala 49:59]
  assign _T_745 = _T_738 ? _T_743 : _T_744; // @[LZD.scala 49:35]
  assign _T_747 = {_T_740,_T_742,_T_745}; // @[Cat.scala 29:58]
  assign _T_748 = _T_686[3]; // @[Shift.scala 12:21]
  assign _T_749 = _T_747[3]; // @[Shift.scala 12:21]
  assign _T_750 = _T_748 | _T_749; // @[LZD.scala 49:16]
  assign _T_751 = ~ _T_749; // @[LZD.scala 49:27]
  assign _T_752 = _T_748 | _T_751; // @[LZD.scala 49:25]
  assign _T_753 = _T_686[2:0]; // @[LZD.scala 49:47]
  assign _T_754 = _T_747[2:0]; // @[LZD.scala 49:59]
  assign _T_755 = _T_748 ? _T_753 : _T_754; // @[LZD.scala 49:35]
  assign _T_757 = {_T_750,_T_752,_T_755}; // @[Cat.scala 29:58]
  assign _T_758 = _T_624[12:0]; // @[LZD.scala 44:32]
  assign _T_759 = _T_758[12:5]; // @[LZD.scala 43:32]
  assign _T_760 = _T_759[7:4]; // @[LZD.scala 43:32]
  assign _T_761 = _T_760[3:2]; // @[LZD.scala 43:32]
  assign _T_762 = _T_761 != 2'h0; // @[LZD.scala 39:14]
  assign _T_763 = _T_761[1]; // @[LZD.scala 39:21]
  assign _T_764 = _T_761[0]; // @[LZD.scala 39:30]
  assign _T_765 = ~ _T_764; // @[LZD.scala 39:27]
  assign _T_766 = _T_763 | _T_765; // @[LZD.scala 39:25]
  assign _T_767 = {_T_762,_T_766}; // @[Cat.scala 29:58]
  assign _T_768 = _T_760[1:0]; // @[LZD.scala 44:32]
  assign _T_769 = _T_768 != 2'h0; // @[LZD.scala 39:14]
  assign _T_770 = _T_768[1]; // @[LZD.scala 39:21]
  assign _T_771 = _T_768[0]; // @[LZD.scala 39:30]
  assign _T_772 = ~ _T_771; // @[LZD.scala 39:27]
  assign _T_773 = _T_770 | _T_772; // @[LZD.scala 39:25]
  assign _T_774 = {_T_769,_T_773}; // @[Cat.scala 29:58]
  assign _T_775 = _T_767[1]; // @[Shift.scala 12:21]
  assign _T_776 = _T_774[1]; // @[Shift.scala 12:21]
  assign _T_777 = _T_775 | _T_776; // @[LZD.scala 49:16]
  assign _T_778 = ~ _T_776; // @[LZD.scala 49:27]
  assign _T_779 = _T_775 | _T_778; // @[LZD.scala 49:25]
  assign _T_780 = _T_767[0:0]; // @[LZD.scala 49:47]
  assign _T_781 = _T_774[0:0]; // @[LZD.scala 49:59]
  assign _T_782 = _T_775 ? _T_780 : _T_781; // @[LZD.scala 49:35]
  assign _T_784 = {_T_777,_T_779,_T_782}; // @[Cat.scala 29:58]
  assign _T_785 = _T_759[3:0]; // @[LZD.scala 44:32]
  assign _T_786 = _T_785[3:2]; // @[LZD.scala 43:32]
  assign _T_787 = _T_786 != 2'h0; // @[LZD.scala 39:14]
  assign _T_788 = _T_786[1]; // @[LZD.scala 39:21]
  assign _T_789 = _T_786[0]; // @[LZD.scala 39:30]
  assign _T_790 = ~ _T_789; // @[LZD.scala 39:27]
  assign _T_791 = _T_788 | _T_790; // @[LZD.scala 39:25]
  assign _T_792 = {_T_787,_T_791}; // @[Cat.scala 29:58]
  assign _T_793 = _T_785[1:0]; // @[LZD.scala 44:32]
  assign _T_794 = _T_793 != 2'h0; // @[LZD.scala 39:14]
  assign _T_795 = _T_793[1]; // @[LZD.scala 39:21]
  assign _T_796 = _T_793[0]; // @[LZD.scala 39:30]
  assign _T_797 = ~ _T_796; // @[LZD.scala 39:27]
  assign _T_798 = _T_795 | _T_797; // @[LZD.scala 39:25]
  assign _T_799 = {_T_794,_T_798}; // @[Cat.scala 29:58]
  assign _T_800 = _T_792[1]; // @[Shift.scala 12:21]
  assign _T_801 = _T_799[1]; // @[Shift.scala 12:21]
  assign _T_802 = _T_800 | _T_801; // @[LZD.scala 49:16]
  assign _T_803 = ~ _T_801; // @[LZD.scala 49:27]
  assign _T_804 = _T_800 | _T_803; // @[LZD.scala 49:25]
  assign _T_805 = _T_792[0:0]; // @[LZD.scala 49:47]
  assign _T_806 = _T_799[0:0]; // @[LZD.scala 49:59]
  assign _T_807 = _T_800 ? _T_805 : _T_806; // @[LZD.scala 49:35]
  assign _T_809 = {_T_802,_T_804,_T_807}; // @[Cat.scala 29:58]
  assign _T_810 = _T_784[2]; // @[Shift.scala 12:21]
  assign _T_811 = _T_809[2]; // @[Shift.scala 12:21]
  assign _T_812 = _T_810 | _T_811; // @[LZD.scala 49:16]
  assign _T_813 = ~ _T_811; // @[LZD.scala 49:27]
  assign _T_814 = _T_810 | _T_813; // @[LZD.scala 49:25]
  assign _T_815 = _T_784[1:0]; // @[LZD.scala 49:47]
  assign _T_816 = _T_809[1:0]; // @[LZD.scala 49:59]
  assign _T_817 = _T_810 ? _T_815 : _T_816; // @[LZD.scala 49:35]
  assign _T_819 = {_T_812,_T_814,_T_817}; // @[Cat.scala 29:58]
  assign _T_820 = _T_758[4:0]; // @[LZD.scala 44:32]
  assign _T_821 = _T_820[4:1]; // @[LZD.scala 43:32]
  assign _T_822 = _T_821[3:2]; // @[LZD.scala 43:32]
  assign _T_823 = _T_822 != 2'h0; // @[LZD.scala 39:14]
  assign _T_824 = _T_822[1]; // @[LZD.scala 39:21]
  assign _T_825 = _T_822[0]; // @[LZD.scala 39:30]
  assign _T_826 = ~ _T_825; // @[LZD.scala 39:27]
  assign _T_827 = _T_824 | _T_826; // @[LZD.scala 39:25]
  assign _T_828 = {_T_823,_T_827}; // @[Cat.scala 29:58]
  assign _T_829 = _T_821[1:0]; // @[LZD.scala 44:32]
  assign _T_830 = _T_829 != 2'h0; // @[LZD.scala 39:14]
  assign _T_831 = _T_829[1]; // @[LZD.scala 39:21]
  assign _T_832 = _T_829[0]; // @[LZD.scala 39:30]
  assign _T_833 = ~ _T_832; // @[LZD.scala 39:27]
  assign _T_834 = _T_831 | _T_833; // @[LZD.scala 39:25]
  assign _T_835 = {_T_830,_T_834}; // @[Cat.scala 29:58]
  assign _T_836 = _T_828[1]; // @[Shift.scala 12:21]
  assign _T_837 = _T_835[1]; // @[Shift.scala 12:21]
  assign _T_838 = _T_836 | _T_837; // @[LZD.scala 49:16]
  assign _T_839 = ~ _T_837; // @[LZD.scala 49:27]
  assign _T_840 = _T_836 | _T_839; // @[LZD.scala 49:25]
  assign _T_841 = _T_828[0:0]; // @[LZD.scala 49:47]
  assign _T_842 = _T_835[0:0]; // @[LZD.scala 49:59]
  assign _T_843 = _T_836 ? _T_841 : _T_842; // @[LZD.scala 49:35]
  assign _T_845 = {_T_838,_T_840,_T_843}; // @[Cat.scala 29:58]
  assign _T_846 = _T_820[0:0]; // @[LZD.scala 44:32]
  assign _T_848 = _T_845[2]; // @[Shift.scala 12:21]
  assign _T_850 = {1'h1,_T_846}; // @[Cat.scala 29:58]
  assign _T_851 = _T_845[1:0]; // @[LZD.scala 55:32]
  assign _T_852 = _T_848 ? _T_851 : _T_850; // @[LZD.scala 55:20]
  assign _T_853 = {_T_848,_T_852}; // @[Cat.scala 29:58]
  assign _T_854 = _T_819[3]; // @[Shift.scala 12:21]
  assign _T_856 = _T_819[2:0]; // @[LZD.scala 55:32]
  assign _T_857 = _T_854 ? _T_856 : _T_853; // @[LZD.scala 55:20]
  assign _T_858 = {_T_854,_T_857}; // @[Cat.scala 29:58]
  assign _T_859 = _T_757[4]; // @[Shift.scala 12:21]
  assign _T_861 = _T_757[3:0]; // @[LZD.scala 55:32]
  assign _T_862 = _T_859 ? _T_861 : _T_858; // @[LZD.scala 55:20]
  assign _T_863 = {_T_859,_T_862}; // @[Cat.scala 29:58]
  assign _T_864 = ~ _T_863; // @[convert.scala 21:22]
  assign _T_865 = realC[27:0]; // @[convert.scala 22:36]
  assign _T_866 = _T_864 < 5'h1c; // @[Shift.scala 16:24]
  assign _T_868 = _T_864[4]; // @[Shift.scala 12:21]
  assign _T_869 = _T_865[11:0]; // @[Shift.scala 64:52]
  assign _T_871 = {_T_869,16'h0}; // @[Cat.scala 29:58]
  assign _T_872 = _T_868 ? _T_871 : _T_865; // @[Shift.scala 64:27]
  assign _T_873 = _T_864[3:0]; // @[Shift.scala 66:70]
  assign _T_874 = _T_873[3]; // @[Shift.scala 12:21]
  assign _T_875 = _T_872[19:0]; // @[Shift.scala 64:52]
  assign _T_877 = {_T_875,8'h0}; // @[Cat.scala 29:58]
  assign _T_878 = _T_874 ? _T_877 : _T_872; // @[Shift.scala 64:27]
  assign _T_879 = _T_873[2:0]; // @[Shift.scala 66:70]
  assign _T_880 = _T_879[2]; // @[Shift.scala 12:21]
  assign _T_881 = _T_878[23:0]; // @[Shift.scala 64:52]
  assign _T_883 = {_T_881,4'h0}; // @[Cat.scala 29:58]
  assign _T_884 = _T_880 ? _T_883 : _T_878; // @[Shift.scala 64:27]
  assign _T_885 = _T_879[1:0]; // @[Shift.scala 66:70]
  assign _T_886 = _T_885[1]; // @[Shift.scala 12:21]
  assign _T_887 = _T_884[25:0]; // @[Shift.scala 64:52]
  assign _T_889 = {_T_887,2'h0}; // @[Cat.scala 29:58]
  assign _T_890 = _T_886 ? _T_889 : _T_884; // @[Shift.scala 64:27]
  assign _T_891 = _T_885[0:0]; // @[Shift.scala 66:70]
  assign _T_893 = _T_890[26:0]; // @[Shift.scala 64:52]
  assign _T_894 = {_T_893,1'h0}; // @[Cat.scala 29:58]
  assign _T_895 = _T_891 ? _T_894 : _T_890; // @[Shift.scala 64:27]
  assign _T_896 = _T_866 ? _T_895 : 28'h0; // @[Shift.scala 16:10]
  assign _T_897 = _T_896[27:25]; // @[convert.scala 23:34]
  assign decC_fraction = _T_896[24:0]; // @[convert.scala 24:34]
  assign _T_899 = _T_621 == 1'h0; // @[convert.scala 25:26]
  assign _T_901 = _T_621 ? _T_864 : _T_863; // @[convert.scala 25:42]
  assign _T_904 = ~ _T_897; // @[convert.scala 26:67]
  assign _T_905 = _T_619 ? _T_904 : _T_897; // @[convert.scala 26:51]
  assign _T_906 = {_T_899,_T_901,_T_905}; // @[Cat.scala 29:58]
  assign _T_908 = realC[29:0]; // @[convert.scala 29:56]
  assign _T_909 = _T_908 != 30'h0; // @[convert.scala 29:60]
  assign _T_910 = ~ _T_909; // @[convert.scala 29:41]
  assign decC_isNaR = _T_619 & _T_910; // @[convert.scala 29:39]
  assign _T_913 = _T_619 == 1'h0; // @[convert.scala 30:19]
  assign decC_isZero = _T_913 & _T_910; // @[convert.scala 30:41]
  assign decC_scale = $signed(_T_906); // @[convert.scala 32:24]
  assign _T_921 = decA_isNaR | decB_isNaR; // @[PositFMA.scala 58:30]
  assign outIsNaR = _T_921 | decC_isNaR; // @[PositFMA.scala 58:44]
  assign _T_922 = ~ _T_13; // @[PositFMA.scala 59:34]
  assign _T_923 = ~ decA_isZero; // @[PositFMA.scala 59:47]
  assign _T_924 = _T_922 & _T_923; // @[PositFMA.scala 59:45]
  assign _T_926 = {_T_13,_T_924,decA_fraction}; // @[Cat.scala 29:58]
  assign sigA = $signed(_T_926); // @[PositFMA.scala 59:76]
  assign _T_927 = ~ _T_316; // @[PositFMA.scala 60:34]
  assign _T_928 = ~ decB_isZero; // @[PositFMA.scala 60:47]
  assign _T_929 = _T_927 & _T_928; // @[PositFMA.scala 60:45]
  assign _T_931 = {_T_316,_T_929,decB_fraction}; // @[Cat.scala 29:58]
  assign sigB = $signed(_T_931); // @[PositFMA.scala 60:76]
  assign _T_932 = $signed(sigA) * $signed(sigB); // @[PositFMA.scala 61:25]
  assign sigP = $unsigned(_T_932); // @[PositFMA.scala 61:33]
  assign head2 = sigP[53:52]; // @[PositFMA.scala 62:28]
  assign _T_933 = head2[1]; // @[PositFMA.scala 63:31]
  assign _T_934 = ~ _T_933; // @[PositFMA.scala 63:25]
  assign _T_935 = head2[0]; // @[PositFMA.scala 63:42]
  assign addTwo = _T_934 & _T_935; // @[PositFMA.scala 63:35]
  assign _T_936 = sigP[53]; // @[PositFMA.scala 65:23]
  assign _T_937 = sigP[51]; // @[PositFMA.scala 65:49]
  assign addOne = _T_936 ^ _T_937; // @[PositFMA.scala 65:43]
  assign _T_938 = {addTwo,addOne}; // @[Cat.scala 29:58]
  assign expBias = {1'b0,$signed(_T_938)}; // @[PositFMA.scala 66:39]
  assign mulSign = sigP[53:53]; // @[PositFMA.scala 67:28]
  assign _T_939 = $signed(decA_scale) + $signed(decB_scale); // @[PositFMA.scala 69:30]
  assign _GEN_12 = {{7{expBias[2]}},expBias}; // @[PositFMA.scala 69:44]
  assign _T_941 = $signed(_T_939) + $signed(_GEN_12); // @[PositFMA.scala 69:44]
  assign mulScale = $signed(_T_941); // @[PositFMA.scala 69:44]
  assign _T_942 = sigP[51:0]; // @[PositFMA.scala 72:29]
  assign _T_943 = sigP[50:0]; // @[PositFMA.scala 73:29]
  assign _T_944 = {_T_943, 1'h0}; // @[PositFMA.scala 73:48]
  assign mulSigTmp = addOne ? _T_942 : _T_944; // @[PositFMA.scala 70:22]
  assign _T_946 = mulSigTmp[51:51]; // @[PositFMA.scala 77:39]
  assign _T_947 = _T_946 | addTwo; // @[PositFMA.scala 77:43]
  assign _T_948 = mulSigTmp[50:0]; // @[PositFMA.scala 78:39]
  assign mulSig = {mulSign,_T_947,_T_948}; // @[Cat.scala 29:58]
  assign _T_974 = ~ addSign_phase2; // @[PositFMA.scala 107:29]
  assign _T_975 = ~ addZero_phase2; // @[PositFMA.scala 107:47]
  assign _T_976 = _T_974 & _T_975; // @[PositFMA.scala 107:45]
  assign extAddSig = {addSign_phase2,_T_976,addFrac_phase2,26'h0}; // @[Cat.scala 29:58]
  assign _GEN_13 = {{1{addScale_phase2[8]}},addScale_phase2}; // @[PositFMA.scala 111:39]
  assign mulGreater = $signed(mulScale_phase2) > $signed(_GEN_13); // @[PositFMA.scala 111:39]
  assign greaterScale = mulGreater ? $signed(mulScale_phase2) : $signed({{1{addScale_phase2[8]}},addScale_phase2}); // @[PositFMA.scala 112:26]
  assign smallerScale = mulGreater ? $signed({{1{addScale_phase2[8]}},addScale_phase2}) : $signed(mulScale_phase2); // @[PositFMA.scala 113:26]
  assign _T_980 = $signed(greaterScale) - $signed(smallerScale); // @[PositFMA.scala 114:36]
  assign scaleDiff = $signed(_T_980); // @[PositFMA.scala 114:36]
  assign greaterSig = mulGreater ? mulSig_phase2 : extAddSig; // @[PositFMA.scala 115:26]
  assign smallerSigTmp = mulGreater ? extAddSig : mulSig_phase2; // @[PositFMA.scala 116:26]
  assign _T_981 = $unsigned(scaleDiff); // @[PositFMA.scala 117:69]
  assign _T_982 = _T_981 < 10'h35; // @[Shift.scala 39:24]
  assign _T_983 = _T_981[5:0]; // @[Shift.scala 40:44]
  assign _T_984 = smallerSigTmp[52:32]; // @[Shift.scala 90:30]
  assign _T_985 = smallerSigTmp[31:0]; // @[Shift.scala 90:48]
  assign _T_986 = _T_985 != 32'h0; // @[Shift.scala 90:57]
  assign _GEN_14 = {{20'd0}, _T_986}; // @[Shift.scala 90:39]
  assign _T_987 = _T_984 | _GEN_14; // @[Shift.scala 90:39]
  assign _T_988 = _T_983[5]; // @[Shift.scala 12:21]
  assign _T_989 = smallerSigTmp[52]; // @[Shift.scala 12:21]
  assign _T_991 = _T_989 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 71:12]
  assign _T_992 = {_T_991,_T_987}; // @[Cat.scala 29:58]
  assign _T_993 = _T_988 ? _T_992 : smallerSigTmp; // @[Shift.scala 91:22]
  assign _T_994 = _T_983[4:0]; // @[Shift.scala 92:77]
  assign _T_995 = _T_993[52:16]; // @[Shift.scala 90:30]
  assign _T_996 = _T_993[15:0]; // @[Shift.scala 90:48]
  assign _T_997 = _T_996 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_15 = {{36'd0}, _T_997}; // @[Shift.scala 90:39]
  assign _T_998 = _T_995 | _GEN_15; // @[Shift.scala 90:39]
  assign _T_999 = _T_994[4]; // @[Shift.scala 12:21]
  assign _T_1000 = _T_993[52]; // @[Shift.scala 12:21]
  assign _T_1002 = _T_1000 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_1003 = {_T_1002,_T_998}; // @[Cat.scala 29:58]
  assign _T_1004 = _T_999 ? _T_1003 : _T_993; // @[Shift.scala 91:22]
  assign _T_1005 = _T_994[3:0]; // @[Shift.scala 92:77]
  assign _T_1006 = _T_1004[52:8]; // @[Shift.scala 90:30]
  assign _T_1007 = _T_1004[7:0]; // @[Shift.scala 90:48]
  assign _T_1008 = _T_1007 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_16 = {{44'd0}, _T_1008}; // @[Shift.scala 90:39]
  assign _T_1009 = _T_1006 | _GEN_16; // @[Shift.scala 90:39]
  assign _T_1010 = _T_1005[3]; // @[Shift.scala 12:21]
  assign _T_1011 = _T_1004[52]; // @[Shift.scala 12:21]
  assign _T_1013 = _T_1011 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_1014 = {_T_1013,_T_1009}; // @[Cat.scala 29:58]
  assign _T_1015 = _T_1010 ? _T_1014 : _T_1004; // @[Shift.scala 91:22]
  assign _T_1016 = _T_1005[2:0]; // @[Shift.scala 92:77]
  assign _T_1017 = _T_1015[52:4]; // @[Shift.scala 90:30]
  assign _T_1018 = _T_1015[3:0]; // @[Shift.scala 90:48]
  assign _T_1019 = _T_1018 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_17 = {{48'd0}, _T_1019}; // @[Shift.scala 90:39]
  assign _T_1020 = _T_1017 | _GEN_17; // @[Shift.scala 90:39]
  assign _T_1021 = _T_1016[2]; // @[Shift.scala 12:21]
  assign _T_1022 = _T_1015[52]; // @[Shift.scala 12:21]
  assign _T_1024 = _T_1022 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_1025 = {_T_1024,_T_1020}; // @[Cat.scala 29:58]
  assign _T_1026 = _T_1021 ? _T_1025 : _T_1015; // @[Shift.scala 91:22]
  assign _T_1027 = _T_1016[1:0]; // @[Shift.scala 92:77]
  assign _T_1028 = _T_1026[52:2]; // @[Shift.scala 90:30]
  assign _T_1029 = _T_1026[1:0]; // @[Shift.scala 90:48]
  assign _T_1030 = _T_1029 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_18 = {{50'd0}, _T_1030}; // @[Shift.scala 90:39]
  assign _T_1031 = _T_1028 | _GEN_18; // @[Shift.scala 90:39]
  assign _T_1032 = _T_1027[1]; // @[Shift.scala 12:21]
  assign _T_1033 = _T_1026[52]; // @[Shift.scala 12:21]
  assign _T_1035 = _T_1033 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_1036 = {_T_1035,_T_1031}; // @[Cat.scala 29:58]
  assign _T_1037 = _T_1032 ? _T_1036 : _T_1026; // @[Shift.scala 91:22]
  assign _T_1038 = _T_1027[0:0]; // @[Shift.scala 92:77]
  assign _T_1039 = _T_1037[52:1]; // @[Shift.scala 90:30]
  assign _T_1040 = _T_1037[0:0]; // @[Shift.scala 90:48]
  assign _GEN_19 = {{51'd0}, _T_1040}; // @[Shift.scala 90:39]
  assign _T_1042 = _T_1039 | _GEN_19; // @[Shift.scala 90:39]
  assign _T_1044 = _T_1037[52]; // @[Shift.scala 12:21]
  assign _T_1045 = {_T_1044,_T_1042}; // @[Cat.scala 29:58]
  assign _T_1046 = _T_1038 ? _T_1045 : _T_1037; // @[Shift.scala 91:22]
  assign _T_1049 = _T_989 ? 53'h1fffffffffffff : 53'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_982 ? _T_1046 : _T_1049; // @[Shift.scala 39:10]
  assign rawSumSig = greaterSig + smallerSig; // @[PositFMA.scala 118:34]
  assign _T_1050 = mulSig_phase2[52:52]; // @[PositFMA.scala 119:42]
  assign _T_1051 = _T_1050 ^ addSign_phase2; // @[PositFMA.scala 119:46]
  assign _T_1052 = rawSumSig[53:53]; // @[PositFMA.scala 119:79]
  assign sumSign = _T_1051 ^ _T_1052; // @[PositFMA.scala 119:63]
  assign _T_1054 = greaterSig + smallerSig; // @[PositFMA.scala 120:50]
  assign signSumSig = {sumSign,_T_1054}; // @[Cat.scala 29:58]
  assign _T_1055 = signSumSig[53:1]; // @[PositFMA.scala 124:33]
  assign _T_1056 = signSumSig[52:0]; // @[PositFMA.scala 124:68]
  assign sumXor = _T_1055 ^ _T_1056; // @[PositFMA.scala 124:51]
  assign _T_1057 = sumXor[52:21]; // @[LZD.scala 43:32]
  assign _T_1058 = _T_1057[31:16]; // @[LZD.scala 43:32]
  assign _T_1059 = _T_1058[15:8]; // @[LZD.scala 43:32]
  assign _T_1060 = _T_1059[7:4]; // @[LZD.scala 43:32]
  assign _T_1061 = _T_1060[3:2]; // @[LZD.scala 43:32]
  assign _T_1062 = _T_1061 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1063 = _T_1061[1]; // @[LZD.scala 39:21]
  assign _T_1064 = _T_1061[0]; // @[LZD.scala 39:30]
  assign _T_1065 = ~ _T_1064; // @[LZD.scala 39:27]
  assign _T_1066 = _T_1063 | _T_1065; // @[LZD.scala 39:25]
  assign _T_1067 = {_T_1062,_T_1066}; // @[Cat.scala 29:58]
  assign _T_1068 = _T_1060[1:0]; // @[LZD.scala 44:32]
  assign _T_1069 = _T_1068 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1070 = _T_1068[1]; // @[LZD.scala 39:21]
  assign _T_1071 = _T_1068[0]; // @[LZD.scala 39:30]
  assign _T_1072 = ~ _T_1071; // @[LZD.scala 39:27]
  assign _T_1073 = _T_1070 | _T_1072; // @[LZD.scala 39:25]
  assign _T_1074 = {_T_1069,_T_1073}; // @[Cat.scala 29:58]
  assign _T_1075 = _T_1067[1]; // @[Shift.scala 12:21]
  assign _T_1076 = _T_1074[1]; // @[Shift.scala 12:21]
  assign _T_1077 = _T_1075 | _T_1076; // @[LZD.scala 49:16]
  assign _T_1078 = ~ _T_1076; // @[LZD.scala 49:27]
  assign _T_1079 = _T_1075 | _T_1078; // @[LZD.scala 49:25]
  assign _T_1080 = _T_1067[0:0]; // @[LZD.scala 49:47]
  assign _T_1081 = _T_1074[0:0]; // @[LZD.scala 49:59]
  assign _T_1082 = _T_1075 ? _T_1080 : _T_1081; // @[LZD.scala 49:35]
  assign _T_1084 = {_T_1077,_T_1079,_T_1082}; // @[Cat.scala 29:58]
  assign _T_1085 = _T_1059[3:0]; // @[LZD.scala 44:32]
  assign _T_1086 = _T_1085[3:2]; // @[LZD.scala 43:32]
  assign _T_1087 = _T_1086 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1088 = _T_1086[1]; // @[LZD.scala 39:21]
  assign _T_1089 = _T_1086[0]; // @[LZD.scala 39:30]
  assign _T_1090 = ~ _T_1089; // @[LZD.scala 39:27]
  assign _T_1091 = _T_1088 | _T_1090; // @[LZD.scala 39:25]
  assign _T_1092 = {_T_1087,_T_1091}; // @[Cat.scala 29:58]
  assign _T_1093 = _T_1085[1:0]; // @[LZD.scala 44:32]
  assign _T_1094 = _T_1093 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1095 = _T_1093[1]; // @[LZD.scala 39:21]
  assign _T_1096 = _T_1093[0]; // @[LZD.scala 39:30]
  assign _T_1097 = ~ _T_1096; // @[LZD.scala 39:27]
  assign _T_1098 = _T_1095 | _T_1097; // @[LZD.scala 39:25]
  assign _T_1099 = {_T_1094,_T_1098}; // @[Cat.scala 29:58]
  assign _T_1100 = _T_1092[1]; // @[Shift.scala 12:21]
  assign _T_1101 = _T_1099[1]; // @[Shift.scala 12:21]
  assign _T_1102 = _T_1100 | _T_1101; // @[LZD.scala 49:16]
  assign _T_1103 = ~ _T_1101; // @[LZD.scala 49:27]
  assign _T_1104 = _T_1100 | _T_1103; // @[LZD.scala 49:25]
  assign _T_1105 = _T_1092[0:0]; // @[LZD.scala 49:47]
  assign _T_1106 = _T_1099[0:0]; // @[LZD.scala 49:59]
  assign _T_1107 = _T_1100 ? _T_1105 : _T_1106; // @[LZD.scala 49:35]
  assign _T_1109 = {_T_1102,_T_1104,_T_1107}; // @[Cat.scala 29:58]
  assign _T_1110 = _T_1084[2]; // @[Shift.scala 12:21]
  assign _T_1111 = _T_1109[2]; // @[Shift.scala 12:21]
  assign _T_1112 = _T_1110 | _T_1111; // @[LZD.scala 49:16]
  assign _T_1113 = ~ _T_1111; // @[LZD.scala 49:27]
  assign _T_1114 = _T_1110 | _T_1113; // @[LZD.scala 49:25]
  assign _T_1115 = _T_1084[1:0]; // @[LZD.scala 49:47]
  assign _T_1116 = _T_1109[1:0]; // @[LZD.scala 49:59]
  assign _T_1117 = _T_1110 ? _T_1115 : _T_1116; // @[LZD.scala 49:35]
  assign _T_1119 = {_T_1112,_T_1114,_T_1117}; // @[Cat.scala 29:58]
  assign _T_1120 = _T_1058[7:0]; // @[LZD.scala 44:32]
  assign _T_1121 = _T_1120[7:4]; // @[LZD.scala 43:32]
  assign _T_1122 = _T_1121[3:2]; // @[LZD.scala 43:32]
  assign _T_1123 = _T_1122 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1124 = _T_1122[1]; // @[LZD.scala 39:21]
  assign _T_1125 = _T_1122[0]; // @[LZD.scala 39:30]
  assign _T_1126 = ~ _T_1125; // @[LZD.scala 39:27]
  assign _T_1127 = _T_1124 | _T_1126; // @[LZD.scala 39:25]
  assign _T_1128 = {_T_1123,_T_1127}; // @[Cat.scala 29:58]
  assign _T_1129 = _T_1121[1:0]; // @[LZD.scala 44:32]
  assign _T_1130 = _T_1129 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1131 = _T_1129[1]; // @[LZD.scala 39:21]
  assign _T_1132 = _T_1129[0]; // @[LZD.scala 39:30]
  assign _T_1133 = ~ _T_1132; // @[LZD.scala 39:27]
  assign _T_1134 = _T_1131 | _T_1133; // @[LZD.scala 39:25]
  assign _T_1135 = {_T_1130,_T_1134}; // @[Cat.scala 29:58]
  assign _T_1136 = _T_1128[1]; // @[Shift.scala 12:21]
  assign _T_1137 = _T_1135[1]; // @[Shift.scala 12:21]
  assign _T_1138 = _T_1136 | _T_1137; // @[LZD.scala 49:16]
  assign _T_1139 = ~ _T_1137; // @[LZD.scala 49:27]
  assign _T_1140 = _T_1136 | _T_1139; // @[LZD.scala 49:25]
  assign _T_1141 = _T_1128[0:0]; // @[LZD.scala 49:47]
  assign _T_1142 = _T_1135[0:0]; // @[LZD.scala 49:59]
  assign _T_1143 = _T_1136 ? _T_1141 : _T_1142; // @[LZD.scala 49:35]
  assign _T_1145 = {_T_1138,_T_1140,_T_1143}; // @[Cat.scala 29:58]
  assign _T_1146 = _T_1120[3:0]; // @[LZD.scala 44:32]
  assign _T_1147 = _T_1146[3:2]; // @[LZD.scala 43:32]
  assign _T_1148 = _T_1147 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1149 = _T_1147[1]; // @[LZD.scala 39:21]
  assign _T_1150 = _T_1147[0]; // @[LZD.scala 39:30]
  assign _T_1151 = ~ _T_1150; // @[LZD.scala 39:27]
  assign _T_1152 = _T_1149 | _T_1151; // @[LZD.scala 39:25]
  assign _T_1153 = {_T_1148,_T_1152}; // @[Cat.scala 29:58]
  assign _T_1154 = _T_1146[1:0]; // @[LZD.scala 44:32]
  assign _T_1155 = _T_1154 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1156 = _T_1154[1]; // @[LZD.scala 39:21]
  assign _T_1157 = _T_1154[0]; // @[LZD.scala 39:30]
  assign _T_1158 = ~ _T_1157; // @[LZD.scala 39:27]
  assign _T_1159 = _T_1156 | _T_1158; // @[LZD.scala 39:25]
  assign _T_1160 = {_T_1155,_T_1159}; // @[Cat.scala 29:58]
  assign _T_1161 = _T_1153[1]; // @[Shift.scala 12:21]
  assign _T_1162 = _T_1160[1]; // @[Shift.scala 12:21]
  assign _T_1163 = _T_1161 | _T_1162; // @[LZD.scala 49:16]
  assign _T_1164 = ~ _T_1162; // @[LZD.scala 49:27]
  assign _T_1165 = _T_1161 | _T_1164; // @[LZD.scala 49:25]
  assign _T_1166 = _T_1153[0:0]; // @[LZD.scala 49:47]
  assign _T_1167 = _T_1160[0:0]; // @[LZD.scala 49:59]
  assign _T_1168 = _T_1161 ? _T_1166 : _T_1167; // @[LZD.scala 49:35]
  assign _T_1170 = {_T_1163,_T_1165,_T_1168}; // @[Cat.scala 29:58]
  assign _T_1171 = _T_1145[2]; // @[Shift.scala 12:21]
  assign _T_1172 = _T_1170[2]; // @[Shift.scala 12:21]
  assign _T_1173 = _T_1171 | _T_1172; // @[LZD.scala 49:16]
  assign _T_1174 = ~ _T_1172; // @[LZD.scala 49:27]
  assign _T_1175 = _T_1171 | _T_1174; // @[LZD.scala 49:25]
  assign _T_1176 = _T_1145[1:0]; // @[LZD.scala 49:47]
  assign _T_1177 = _T_1170[1:0]; // @[LZD.scala 49:59]
  assign _T_1178 = _T_1171 ? _T_1176 : _T_1177; // @[LZD.scala 49:35]
  assign _T_1180 = {_T_1173,_T_1175,_T_1178}; // @[Cat.scala 29:58]
  assign _T_1181 = _T_1119[3]; // @[Shift.scala 12:21]
  assign _T_1182 = _T_1180[3]; // @[Shift.scala 12:21]
  assign _T_1183 = _T_1181 | _T_1182; // @[LZD.scala 49:16]
  assign _T_1184 = ~ _T_1182; // @[LZD.scala 49:27]
  assign _T_1185 = _T_1181 | _T_1184; // @[LZD.scala 49:25]
  assign _T_1186 = _T_1119[2:0]; // @[LZD.scala 49:47]
  assign _T_1187 = _T_1180[2:0]; // @[LZD.scala 49:59]
  assign _T_1188 = _T_1181 ? _T_1186 : _T_1187; // @[LZD.scala 49:35]
  assign _T_1190 = {_T_1183,_T_1185,_T_1188}; // @[Cat.scala 29:58]
  assign _T_1191 = _T_1057[15:0]; // @[LZD.scala 44:32]
  assign _T_1192 = _T_1191[15:8]; // @[LZD.scala 43:32]
  assign _T_1193 = _T_1192[7:4]; // @[LZD.scala 43:32]
  assign _T_1194 = _T_1193[3:2]; // @[LZD.scala 43:32]
  assign _T_1195 = _T_1194 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1196 = _T_1194[1]; // @[LZD.scala 39:21]
  assign _T_1197 = _T_1194[0]; // @[LZD.scala 39:30]
  assign _T_1198 = ~ _T_1197; // @[LZD.scala 39:27]
  assign _T_1199 = _T_1196 | _T_1198; // @[LZD.scala 39:25]
  assign _T_1200 = {_T_1195,_T_1199}; // @[Cat.scala 29:58]
  assign _T_1201 = _T_1193[1:0]; // @[LZD.scala 44:32]
  assign _T_1202 = _T_1201 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1203 = _T_1201[1]; // @[LZD.scala 39:21]
  assign _T_1204 = _T_1201[0]; // @[LZD.scala 39:30]
  assign _T_1205 = ~ _T_1204; // @[LZD.scala 39:27]
  assign _T_1206 = _T_1203 | _T_1205; // @[LZD.scala 39:25]
  assign _T_1207 = {_T_1202,_T_1206}; // @[Cat.scala 29:58]
  assign _T_1208 = _T_1200[1]; // @[Shift.scala 12:21]
  assign _T_1209 = _T_1207[1]; // @[Shift.scala 12:21]
  assign _T_1210 = _T_1208 | _T_1209; // @[LZD.scala 49:16]
  assign _T_1211 = ~ _T_1209; // @[LZD.scala 49:27]
  assign _T_1212 = _T_1208 | _T_1211; // @[LZD.scala 49:25]
  assign _T_1213 = _T_1200[0:0]; // @[LZD.scala 49:47]
  assign _T_1214 = _T_1207[0:0]; // @[LZD.scala 49:59]
  assign _T_1215 = _T_1208 ? _T_1213 : _T_1214; // @[LZD.scala 49:35]
  assign _T_1217 = {_T_1210,_T_1212,_T_1215}; // @[Cat.scala 29:58]
  assign _T_1218 = _T_1192[3:0]; // @[LZD.scala 44:32]
  assign _T_1219 = _T_1218[3:2]; // @[LZD.scala 43:32]
  assign _T_1220 = _T_1219 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1221 = _T_1219[1]; // @[LZD.scala 39:21]
  assign _T_1222 = _T_1219[0]; // @[LZD.scala 39:30]
  assign _T_1223 = ~ _T_1222; // @[LZD.scala 39:27]
  assign _T_1224 = _T_1221 | _T_1223; // @[LZD.scala 39:25]
  assign _T_1225 = {_T_1220,_T_1224}; // @[Cat.scala 29:58]
  assign _T_1226 = _T_1218[1:0]; // @[LZD.scala 44:32]
  assign _T_1227 = _T_1226 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1228 = _T_1226[1]; // @[LZD.scala 39:21]
  assign _T_1229 = _T_1226[0]; // @[LZD.scala 39:30]
  assign _T_1230 = ~ _T_1229; // @[LZD.scala 39:27]
  assign _T_1231 = _T_1228 | _T_1230; // @[LZD.scala 39:25]
  assign _T_1232 = {_T_1227,_T_1231}; // @[Cat.scala 29:58]
  assign _T_1233 = _T_1225[1]; // @[Shift.scala 12:21]
  assign _T_1234 = _T_1232[1]; // @[Shift.scala 12:21]
  assign _T_1235 = _T_1233 | _T_1234; // @[LZD.scala 49:16]
  assign _T_1236 = ~ _T_1234; // @[LZD.scala 49:27]
  assign _T_1237 = _T_1233 | _T_1236; // @[LZD.scala 49:25]
  assign _T_1238 = _T_1225[0:0]; // @[LZD.scala 49:47]
  assign _T_1239 = _T_1232[0:0]; // @[LZD.scala 49:59]
  assign _T_1240 = _T_1233 ? _T_1238 : _T_1239; // @[LZD.scala 49:35]
  assign _T_1242 = {_T_1235,_T_1237,_T_1240}; // @[Cat.scala 29:58]
  assign _T_1243 = _T_1217[2]; // @[Shift.scala 12:21]
  assign _T_1244 = _T_1242[2]; // @[Shift.scala 12:21]
  assign _T_1245 = _T_1243 | _T_1244; // @[LZD.scala 49:16]
  assign _T_1246 = ~ _T_1244; // @[LZD.scala 49:27]
  assign _T_1247 = _T_1243 | _T_1246; // @[LZD.scala 49:25]
  assign _T_1248 = _T_1217[1:0]; // @[LZD.scala 49:47]
  assign _T_1249 = _T_1242[1:0]; // @[LZD.scala 49:59]
  assign _T_1250 = _T_1243 ? _T_1248 : _T_1249; // @[LZD.scala 49:35]
  assign _T_1252 = {_T_1245,_T_1247,_T_1250}; // @[Cat.scala 29:58]
  assign _T_1253 = _T_1191[7:0]; // @[LZD.scala 44:32]
  assign _T_1254 = _T_1253[7:4]; // @[LZD.scala 43:32]
  assign _T_1255 = _T_1254[3:2]; // @[LZD.scala 43:32]
  assign _T_1256 = _T_1255 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1257 = _T_1255[1]; // @[LZD.scala 39:21]
  assign _T_1258 = _T_1255[0]; // @[LZD.scala 39:30]
  assign _T_1259 = ~ _T_1258; // @[LZD.scala 39:27]
  assign _T_1260 = _T_1257 | _T_1259; // @[LZD.scala 39:25]
  assign _T_1261 = {_T_1256,_T_1260}; // @[Cat.scala 29:58]
  assign _T_1262 = _T_1254[1:0]; // @[LZD.scala 44:32]
  assign _T_1263 = _T_1262 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1264 = _T_1262[1]; // @[LZD.scala 39:21]
  assign _T_1265 = _T_1262[0]; // @[LZD.scala 39:30]
  assign _T_1266 = ~ _T_1265; // @[LZD.scala 39:27]
  assign _T_1267 = _T_1264 | _T_1266; // @[LZD.scala 39:25]
  assign _T_1268 = {_T_1263,_T_1267}; // @[Cat.scala 29:58]
  assign _T_1269 = _T_1261[1]; // @[Shift.scala 12:21]
  assign _T_1270 = _T_1268[1]; // @[Shift.scala 12:21]
  assign _T_1271 = _T_1269 | _T_1270; // @[LZD.scala 49:16]
  assign _T_1272 = ~ _T_1270; // @[LZD.scala 49:27]
  assign _T_1273 = _T_1269 | _T_1272; // @[LZD.scala 49:25]
  assign _T_1274 = _T_1261[0:0]; // @[LZD.scala 49:47]
  assign _T_1275 = _T_1268[0:0]; // @[LZD.scala 49:59]
  assign _T_1276 = _T_1269 ? _T_1274 : _T_1275; // @[LZD.scala 49:35]
  assign _T_1278 = {_T_1271,_T_1273,_T_1276}; // @[Cat.scala 29:58]
  assign _T_1279 = _T_1253[3:0]; // @[LZD.scala 44:32]
  assign _T_1280 = _T_1279[3:2]; // @[LZD.scala 43:32]
  assign _T_1281 = _T_1280 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1282 = _T_1280[1]; // @[LZD.scala 39:21]
  assign _T_1283 = _T_1280[0]; // @[LZD.scala 39:30]
  assign _T_1284 = ~ _T_1283; // @[LZD.scala 39:27]
  assign _T_1285 = _T_1282 | _T_1284; // @[LZD.scala 39:25]
  assign _T_1286 = {_T_1281,_T_1285}; // @[Cat.scala 29:58]
  assign _T_1287 = _T_1279[1:0]; // @[LZD.scala 44:32]
  assign _T_1288 = _T_1287 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1289 = _T_1287[1]; // @[LZD.scala 39:21]
  assign _T_1290 = _T_1287[0]; // @[LZD.scala 39:30]
  assign _T_1291 = ~ _T_1290; // @[LZD.scala 39:27]
  assign _T_1292 = _T_1289 | _T_1291; // @[LZD.scala 39:25]
  assign _T_1293 = {_T_1288,_T_1292}; // @[Cat.scala 29:58]
  assign _T_1294 = _T_1286[1]; // @[Shift.scala 12:21]
  assign _T_1295 = _T_1293[1]; // @[Shift.scala 12:21]
  assign _T_1296 = _T_1294 | _T_1295; // @[LZD.scala 49:16]
  assign _T_1297 = ~ _T_1295; // @[LZD.scala 49:27]
  assign _T_1298 = _T_1294 | _T_1297; // @[LZD.scala 49:25]
  assign _T_1299 = _T_1286[0:0]; // @[LZD.scala 49:47]
  assign _T_1300 = _T_1293[0:0]; // @[LZD.scala 49:59]
  assign _T_1301 = _T_1294 ? _T_1299 : _T_1300; // @[LZD.scala 49:35]
  assign _T_1303 = {_T_1296,_T_1298,_T_1301}; // @[Cat.scala 29:58]
  assign _T_1304 = _T_1278[2]; // @[Shift.scala 12:21]
  assign _T_1305 = _T_1303[2]; // @[Shift.scala 12:21]
  assign _T_1306 = _T_1304 | _T_1305; // @[LZD.scala 49:16]
  assign _T_1307 = ~ _T_1305; // @[LZD.scala 49:27]
  assign _T_1308 = _T_1304 | _T_1307; // @[LZD.scala 49:25]
  assign _T_1309 = _T_1278[1:0]; // @[LZD.scala 49:47]
  assign _T_1310 = _T_1303[1:0]; // @[LZD.scala 49:59]
  assign _T_1311 = _T_1304 ? _T_1309 : _T_1310; // @[LZD.scala 49:35]
  assign _T_1313 = {_T_1306,_T_1308,_T_1311}; // @[Cat.scala 29:58]
  assign _T_1314 = _T_1252[3]; // @[Shift.scala 12:21]
  assign _T_1315 = _T_1313[3]; // @[Shift.scala 12:21]
  assign _T_1316 = _T_1314 | _T_1315; // @[LZD.scala 49:16]
  assign _T_1317 = ~ _T_1315; // @[LZD.scala 49:27]
  assign _T_1318 = _T_1314 | _T_1317; // @[LZD.scala 49:25]
  assign _T_1319 = _T_1252[2:0]; // @[LZD.scala 49:47]
  assign _T_1320 = _T_1313[2:0]; // @[LZD.scala 49:59]
  assign _T_1321 = _T_1314 ? _T_1319 : _T_1320; // @[LZD.scala 49:35]
  assign _T_1323 = {_T_1316,_T_1318,_T_1321}; // @[Cat.scala 29:58]
  assign _T_1324 = _T_1190[4]; // @[Shift.scala 12:21]
  assign _T_1325 = _T_1323[4]; // @[Shift.scala 12:21]
  assign _T_1326 = _T_1324 | _T_1325; // @[LZD.scala 49:16]
  assign _T_1327 = ~ _T_1325; // @[LZD.scala 49:27]
  assign _T_1328 = _T_1324 | _T_1327; // @[LZD.scala 49:25]
  assign _T_1329 = _T_1190[3:0]; // @[LZD.scala 49:47]
  assign _T_1330 = _T_1323[3:0]; // @[LZD.scala 49:59]
  assign _T_1331 = _T_1324 ? _T_1329 : _T_1330; // @[LZD.scala 49:35]
  assign _T_1333 = {_T_1326,_T_1328,_T_1331}; // @[Cat.scala 29:58]
  assign _T_1334 = sumXor[20:0]; // @[LZD.scala 44:32]
  assign _T_1335 = _T_1334[20:5]; // @[LZD.scala 43:32]
  assign _T_1336 = _T_1335[15:8]; // @[LZD.scala 43:32]
  assign _T_1337 = _T_1336[7:4]; // @[LZD.scala 43:32]
  assign _T_1338 = _T_1337[3:2]; // @[LZD.scala 43:32]
  assign _T_1339 = _T_1338 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1340 = _T_1338[1]; // @[LZD.scala 39:21]
  assign _T_1341 = _T_1338[0]; // @[LZD.scala 39:30]
  assign _T_1342 = ~ _T_1341; // @[LZD.scala 39:27]
  assign _T_1343 = _T_1340 | _T_1342; // @[LZD.scala 39:25]
  assign _T_1344 = {_T_1339,_T_1343}; // @[Cat.scala 29:58]
  assign _T_1345 = _T_1337[1:0]; // @[LZD.scala 44:32]
  assign _T_1346 = _T_1345 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1347 = _T_1345[1]; // @[LZD.scala 39:21]
  assign _T_1348 = _T_1345[0]; // @[LZD.scala 39:30]
  assign _T_1349 = ~ _T_1348; // @[LZD.scala 39:27]
  assign _T_1350 = _T_1347 | _T_1349; // @[LZD.scala 39:25]
  assign _T_1351 = {_T_1346,_T_1350}; // @[Cat.scala 29:58]
  assign _T_1352 = _T_1344[1]; // @[Shift.scala 12:21]
  assign _T_1353 = _T_1351[1]; // @[Shift.scala 12:21]
  assign _T_1354 = _T_1352 | _T_1353; // @[LZD.scala 49:16]
  assign _T_1355 = ~ _T_1353; // @[LZD.scala 49:27]
  assign _T_1356 = _T_1352 | _T_1355; // @[LZD.scala 49:25]
  assign _T_1357 = _T_1344[0:0]; // @[LZD.scala 49:47]
  assign _T_1358 = _T_1351[0:0]; // @[LZD.scala 49:59]
  assign _T_1359 = _T_1352 ? _T_1357 : _T_1358; // @[LZD.scala 49:35]
  assign _T_1361 = {_T_1354,_T_1356,_T_1359}; // @[Cat.scala 29:58]
  assign _T_1362 = _T_1336[3:0]; // @[LZD.scala 44:32]
  assign _T_1363 = _T_1362[3:2]; // @[LZD.scala 43:32]
  assign _T_1364 = _T_1363 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1365 = _T_1363[1]; // @[LZD.scala 39:21]
  assign _T_1366 = _T_1363[0]; // @[LZD.scala 39:30]
  assign _T_1367 = ~ _T_1366; // @[LZD.scala 39:27]
  assign _T_1368 = _T_1365 | _T_1367; // @[LZD.scala 39:25]
  assign _T_1369 = {_T_1364,_T_1368}; // @[Cat.scala 29:58]
  assign _T_1370 = _T_1362[1:0]; // @[LZD.scala 44:32]
  assign _T_1371 = _T_1370 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1372 = _T_1370[1]; // @[LZD.scala 39:21]
  assign _T_1373 = _T_1370[0]; // @[LZD.scala 39:30]
  assign _T_1374 = ~ _T_1373; // @[LZD.scala 39:27]
  assign _T_1375 = _T_1372 | _T_1374; // @[LZD.scala 39:25]
  assign _T_1376 = {_T_1371,_T_1375}; // @[Cat.scala 29:58]
  assign _T_1377 = _T_1369[1]; // @[Shift.scala 12:21]
  assign _T_1378 = _T_1376[1]; // @[Shift.scala 12:21]
  assign _T_1379 = _T_1377 | _T_1378; // @[LZD.scala 49:16]
  assign _T_1380 = ~ _T_1378; // @[LZD.scala 49:27]
  assign _T_1381 = _T_1377 | _T_1380; // @[LZD.scala 49:25]
  assign _T_1382 = _T_1369[0:0]; // @[LZD.scala 49:47]
  assign _T_1383 = _T_1376[0:0]; // @[LZD.scala 49:59]
  assign _T_1384 = _T_1377 ? _T_1382 : _T_1383; // @[LZD.scala 49:35]
  assign _T_1386 = {_T_1379,_T_1381,_T_1384}; // @[Cat.scala 29:58]
  assign _T_1387 = _T_1361[2]; // @[Shift.scala 12:21]
  assign _T_1388 = _T_1386[2]; // @[Shift.scala 12:21]
  assign _T_1389 = _T_1387 | _T_1388; // @[LZD.scala 49:16]
  assign _T_1390 = ~ _T_1388; // @[LZD.scala 49:27]
  assign _T_1391 = _T_1387 | _T_1390; // @[LZD.scala 49:25]
  assign _T_1392 = _T_1361[1:0]; // @[LZD.scala 49:47]
  assign _T_1393 = _T_1386[1:0]; // @[LZD.scala 49:59]
  assign _T_1394 = _T_1387 ? _T_1392 : _T_1393; // @[LZD.scala 49:35]
  assign _T_1396 = {_T_1389,_T_1391,_T_1394}; // @[Cat.scala 29:58]
  assign _T_1397 = _T_1335[7:0]; // @[LZD.scala 44:32]
  assign _T_1398 = _T_1397[7:4]; // @[LZD.scala 43:32]
  assign _T_1399 = _T_1398[3:2]; // @[LZD.scala 43:32]
  assign _T_1400 = _T_1399 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1401 = _T_1399[1]; // @[LZD.scala 39:21]
  assign _T_1402 = _T_1399[0]; // @[LZD.scala 39:30]
  assign _T_1403 = ~ _T_1402; // @[LZD.scala 39:27]
  assign _T_1404 = _T_1401 | _T_1403; // @[LZD.scala 39:25]
  assign _T_1405 = {_T_1400,_T_1404}; // @[Cat.scala 29:58]
  assign _T_1406 = _T_1398[1:0]; // @[LZD.scala 44:32]
  assign _T_1407 = _T_1406 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1408 = _T_1406[1]; // @[LZD.scala 39:21]
  assign _T_1409 = _T_1406[0]; // @[LZD.scala 39:30]
  assign _T_1410 = ~ _T_1409; // @[LZD.scala 39:27]
  assign _T_1411 = _T_1408 | _T_1410; // @[LZD.scala 39:25]
  assign _T_1412 = {_T_1407,_T_1411}; // @[Cat.scala 29:58]
  assign _T_1413 = _T_1405[1]; // @[Shift.scala 12:21]
  assign _T_1414 = _T_1412[1]; // @[Shift.scala 12:21]
  assign _T_1415 = _T_1413 | _T_1414; // @[LZD.scala 49:16]
  assign _T_1416 = ~ _T_1414; // @[LZD.scala 49:27]
  assign _T_1417 = _T_1413 | _T_1416; // @[LZD.scala 49:25]
  assign _T_1418 = _T_1405[0:0]; // @[LZD.scala 49:47]
  assign _T_1419 = _T_1412[0:0]; // @[LZD.scala 49:59]
  assign _T_1420 = _T_1413 ? _T_1418 : _T_1419; // @[LZD.scala 49:35]
  assign _T_1422 = {_T_1415,_T_1417,_T_1420}; // @[Cat.scala 29:58]
  assign _T_1423 = _T_1397[3:0]; // @[LZD.scala 44:32]
  assign _T_1424 = _T_1423[3:2]; // @[LZD.scala 43:32]
  assign _T_1425 = _T_1424 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1426 = _T_1424[1]; // @[LZD.scala 39:21]
  assign _T_1427 = _T_1424[0]; // @[LZD.scala 39:30]
  assign _T_1428 = ~ _T_1427; // @[LZD.scala 39:27]
  assign _T_1429 = _T_1426 | _T_1428; // @[LZD.scala 39:25]
  assign _T_1430 = {_T_1425,_T_1429}; // @[Cat.scala 29:58]
  assign _T_1431 = _T_1423[1:0]; // @[LZD.scala 44:32]
  assign _T_1432 = _T_1431 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1433 = _T_1431[1]; // @[LZD.scala 39:21]
  assign _T_1434 = _T_1431[0]; // @[LZD.scala 39:30]
  assign _T_1435 = ~ _T_1434; // @[LZD.scala 39:27]
  assign _T_1436 = _T_1433 | _T_1435; // @[LZD.scala 39:25]
  assign _T_1437 = {_T_1432,_T_1436}; // @[Cat.scala 29:58]
  assign _T_1438 = _T_1430[1]; // @[Shift.scala 12:21]
  assign _T_1439 = _T_1437[1]; // @[Shift.scala 12:21]
  assign _T_1440 = _T_1438 | _T_1439; // @[LZD.scala 49:16]
  assign _T_1441 = ~ _T_1439; // @[LZD.scala 49:27]
  assign _T_1442 = _T_1438 | _T_1441; // @[LZD.scala 49:25]
  assign _T_1443 = _T_1430[0:0]; // @[LZD.scala 49:47]
  assign _T_1444 = _T_1437[0:0]; // @[LZD.scala 49:59]
  assign _T_1445 = _T_1438 ? _T_1443 : _T_1444; // @[LZD.scala 49:35]
  assign _T_1447 = {_T_1440,_T_1442,_T_1445}; // @[Cat.scala 29:58]
  assign _T_1448 = _T_1422[2]; // @[Shift.scala 12:21]
  assign _T_1449 = _T_1447[2]; // @[Shift.scala 12:21]
  assign _T_1450 = _T_1448 | _T_1449; // @[LZD.scala 49:16]
  assign _T_1451 = ~ _T_1449; // @[LZD.scala 49:27]
  assign _T_1452 = _T_1448 | _T_1451; // @[LZD.scala 49:25]
  assign _T_1453 = _T_1422[1:0]; // @[LZD.scala 49:47]
  assign _T_1454 = _T_1447[1:0]; // @[LZD.scala 49:59]
  assign _T_1455 = _T_1448 ? _T_1453 : _T_1454; // @[LZD.scala 49:35]
  assign _T_1457 = {_T_1450,_T_1452,_T_1455}; // @[Cat.scala 29:58]
  assign _T_1458 = _T_1396[3]; // @[Shift.scala 12:21]
  assign _T_1459 = _T_1457[3]; // @[Shift.scala 12:21]
  assign _T_1460 = _T_1458 | _T_1459; // @[LZD.scala 49:16]
  assign _T_1461 = ~ _T_1459; // @[LZD.scala 49:27]
  assign _T_1462 = _T_1458 | _T_1461; // @[LZD.scala 49:25]
  assign _T_1463 = _T_1396[2:0]; // @[LZD.scala 49:47]
  assign _T_1464 = _T_1457[2:0]; // @[LZD.scala 49:59]
  assign _T_1465 = _T_1458 ? _T_1463 : _T_1464; // @[LZD.scala 49:35]
  assign _T_1467 = {_T_1460,_T_1462,_T_1465}; // @[Cat.scala 29:58]
  assign _T_1468 = _T_1334[4:0]; // @[LZD.scala 44:32]
  assign _T_1469 = _T_1468[4:1]; // @[LZD.scala 43:32]
  assign _T_1470 = _T_1469[3:2]; // @[LZD.scala 43:32]
  assign _T_1471 = _T_1470 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1472 = _T_1470[1]; // @[LZD.scala 39:21]
  assign _T_1473 = _T_1470[0]; // @[LZD.scala 39:30]
  assign _T_1474 = ~ _T_1473; // @[LZD.scala 39:27]
  assign _T_1475 = _T_1472 | _T_1474; // @[LZD.scala 39:25]
  assign _T_1476 = {_T_1471,_T_1475}; // @[Cat.scala 29:58]
  assign _T_1477 = _T_1469[1:0]; // @[LZD.scala 44:32]
  assign _T_1478 = _T_1477 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1479 = _T_1477[1]; // @[LZD.scala 39:21]
  assign _T_1480 = _T_1477[0]; // @[LZD.scala 39:30]
  assign _T_1481 = ~ _T_1480; // @[LZD.scala 39:27]
  assign _T_1482 = _T_1479 | _T_1481; // @[LZD.scala 39:25]
  assign _T_1483 = {_T_1478,_T_1482}; // @[Cat.scala 29:58]
  assign _T_1484 = _T_1476[1]; // @[Shift.scala 12:21]
  assign _T_1485 = _T_1483[1]; // @[Shift.scala 12:21]
  assign _T_1486 = _T_1484 | _T_1485; // @[LZD.scala 49:16]
  assign _T_1487 = ~ _T_1485; // @[LZD.scala 49:27]
  assign _T_1488 = _T_1484 | _T_1487; // @[LZD.scala 49:25]
  assign _T_1489 = _T_1476[0:0]; // @[LZD.scala 49:47]
  assign _T_1490 = _T_1483[0:0]; // @[LZD.scala 49:59]
  assign _T_1491 = _T_1484 ? _T_1489 : _T_1490; // @[LZD.scala 49:35]
  assign _T_1493 = {_T_1486,_T_1488,_T_1491}; // @[Cat.scala 29:58]
  assign _T_1494 = _T_1468[0:0]; // @[LZD.scala 44:32]
  assign _T_1496 = _T_1493[2]; // @[Shift.scala 12:21]
  assign _T_1498 = {1'h1,_T_1494}; // @[Cat.scala 29:58]
  assign _T_1499 = _T_1493[1:0]; // @[LZD.scala 55:32]
  assign _T_1500 = _T_1496 ? _T_1499 : _T_1498; // @[LZD.scala 55:20]
  assign _T_1502 = _T_1467[4]; // @[Shift.scala 12:21]
  assign _T_1504 = {1'h1,_T_1496,_T_1500}; // @[Cat.scala 29:58]
  assign _T_1505 = _T_1467[3:0]; // @[LZD.scala 55:32]
  assign _T_1506 = _T_1502 ? _T_1505 : _T_1504; // @[LZD.scala 55:20]
  assign _T_1507 = {_T_1502,_T_1506}; // @[Cat.scala 29:58]
  assign _T_1508 = _T_1333[5]; // @[Shift.scala 12:21]
  assign _T_1510 = _T_1333[4:0]; // @[LZD.scala 55:32]
  assign _T_1511 = _T_1508 ? _T_1510 : _T_1507; // @[LZD.scala 55:20]
  assign sumLZD = {_T_1508,_T_1511}; // @[Cat.scala 29:58]
  assign shiftValue = ~ sumLZD; // @[PositFMA.scala 126:24]
  assign _T_1512 = signSumSig[51:0]; // @[PositFMA.scala 127:38]
  assign _T_1513 = shiftValue < 6'h34; // @[Shift.scala 16:24]
  assign _T_1515 = shiftValue[5]; // @[Shift.scala 12:21]
  assign _T_1516 = _T_1512[19:0]; // @[Shift.scala 64:52]
  assign _T_1518 = {_T_1516,32'h0}; // @[Cat.scala 29:58]
  assign _T_1519 = _T_1515 ? _T_1518 : _T_1512; // @[Shift.scala 64:27]
  assign _T_1520 = shiftValue[4:0]; // @[Shift.scala 66:70]
  assign _T_1521 = _T_1520[4]; // @[Shift.scala 12:21]
  assign _T_1522 = _T_1519[35:0]; // @[Shift.scala 64:52]
  assign _T_1524 = {_T_1522,16'h0}; // @[Cat.scala 29:58]
  assign _T_1525 = _T_1521 ? _T_1524 : _T_1519; // @[Shift.scala 64:27]
  assign _T_1526 = _T_1520[3:0]; // @[Shift.scala 66:70]
  assign _T_1527 = _T_1526[3]; // @[Shift.scala 12:21]
  assign _T_1528 = _T_1525[43:0]; // @[Shift.scala 64:52]
  assign _T_1530 = {_T_1528,8'h0}; // @[Cat.scala 29:58]
  assign _T_1531 = _T_1527 ? _T_1530 : _T_1525; // @[Shift.scala 64:27]
  assign _T_1532 = _T_1526[2:0]; // @[Shift.scala 66:70]
  assign _T_1533 = _T_1532[2]; // @[Shift.scala 12:21]
  assign _T_1534 = _T_1531[47:0]; // @[Shift.scala 64:52]
  assign _T_1536 = {_T_1534,4'h0}; // @[Cat.scala 29:58]
  assign _T_1537 = _T_1533 ? _T_1536 : _T_1531; // @[Shift.scala 64:27]
  assign _T_1538 = _T_1532[1:0]; // @[Shift.scala 66:70]
  assign _T_1539 = _T_1538[1]; // @[Shift.scala 12:21]
  assign _T_1540 = _T_1537[49:0]; // @[Shift.scala 64:52]
  assign _T_1542 = {_T_1540,2'h0}; // @[Cat.scala 29:58]
  assign _T_1543 = _T_1539 ? _T_1542 : _T_1537; // @[Shift.scala 64:27]
  assign _T_1544 = _T_1538[0:0]; // @[Shift.scala 66:70]
  assign _T_1546 = _T_1543[50:0]; // @[Shift.scala 64:52]
  assign _T_1547 = {_T_1546,1'h0}; // @[Cat.scala 29:58]
  assign _T_1548 = _T_1544 ? _T_1547 : _T_1543; // @[Shift.scala 64:27]
  assign normalFracTmp = _T_1513 ? _T_1548 : 52'h0; // @[Shift.scala 16:10]
  assign _T_1550 = $signed(greaterScale) + $signed(10'sh2); // @[PositFMA.scala 130:36]
  assign _T_1551 = $signed(_T_1550); // @[PositFMA.scala 130:36]
  assign _T_1552 = {1'h1,_T_1508,_T_1511}; // @[Cat.scala 29:58]
  assign _T_1553 = $signed(_T_1552); // @[PositFMA.scala 130:61]
  assign _GEN_20 = {{3{_T_1553[6]}},_T_1553}; // @[PositFMA.scala 130:42]
  assign _T_1555 = $signed(_T_1551) + $signed(_GEN_20); // @[PositFMA.scala 130:42]
  assign sumScale = $signed(_T_1555); // @[PositFMA.scala 130:42]
  assign sumFrac = normalFracTmp[51:27]; // @[PositFMA.scala 131:41]
  assign grsTmp = normalFracTmp[26:0]; // @[PositFMA.scala 134:41]
  assign _T_1556 = grsTmp[26:25]; // @[PositFMA.scala 137:40]
  assign _T_1557 = grsTmp[24:0]; // @[PositFMA.scala 137:56]
  assign _T_1558 = _T_1557 != 25'h0; // @[PositFMA.scala 137:60]
  assign underflow = $signed(sumScale) < $signed(-10'she9); // @[PositFMA.scala 144:32]
  assign overflow = $signed(sumScale) > $signed(10'she8); // @[PositFMA.scala 145:32]
  assign _T_1559 = signSumSig != 54'h0; // @[PositFMA.scala 154:32]
  assign decF_isZero = ~ _T_1559; // @[PositFMA.scala 154:20]
  assign _T_1561 = underflow ? $signed(-10'she9) : $signed(sumScale); // @[Mux.scala 87:16]
  assign _T_1562 = overflow ? $signed(10'she8) : $signed(_T_1561); // @[Mux.scala 87:16]
  assign _GEN_21 = _T_1562[8:0]; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  assign decF_scale = $signed(_GEN_21); // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  assign _T_1563 = decF_scale[2:0]; // @[convert.scala 46:61]
  assign _T_1564 = ~ _T_1563; // @[convert.scala 46:52]
  assign _T_1566 = sumSign ? _T_1564 : _T_1563; // @[convert.scala 46:42]
  assign _T_1567 = decF_scale[8:3]; // @[convert.scala 48:34]
  assign _T_1568 = _T_1567[5:5]; // @[convert.scala 49:36]
  assign _T_1570 = ~ _T_1567; // @[convert.scala 50:36]
  assign _T_1571 = $signed(_T_1570); // @[convert.scala 50:36]
  assign _T_1572 = _T_1568 ? $signed(_T_1571) : $signed(_T_1567); // @[convert.scala 50:28]
  assign _T_1573 = _T_1568 ^ sumSign; // @[convert.scala 51:31]
  assign _T_1574 = ~ _T_1573; // @[convert.scala 52:43]
  assign _T_1578 = {_T_1574,_T_1573,_T_1566,sumFrac,_T_1556,_T_1558}; // @[Cat.scala 29:58]
  assign _T_1579 = $unsigned(_T_1572); // @[Shift.scala 39:17]
  assign _T_1580 = _T_1579 < 6'h21; // @[Shift.scala 39:24]
  assign _T_1582 = _T_1578[32:32]; // @[Shift.scala 90:30]
  assign _T_1583 = _T_1578[31:0]; // @[Shift.scala 90:48]
  assign _T_1584 = _T_1583 != 32'h0; // @[Shift.scala 90:57]
  assign _T_1585 = _T_1582 | _T_1584; // @[Shift.scala 90:39]
  assign _T_1586 = _T_1579[5]; // @[Shift.scala 12:21]
  assign _T_1587 = _T_1578[32]; // @[Shift.scala 12:21]
  assign _T_1589 = _T_1587 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 71:12]
  assign _T_1590 = {_T_1589,_T_1585}; // @[Cat.scala 29:58]
  assign _T_1591 = _T_1586 ? _T_1590 : _T_1578; // @[Shift.scala 91:22]
  assign _T_1592 = _T_1579[4:0]; // @[Shift.scala 92:77]
  assign _T_1593 = _T_1591[32:16]; // @[Shift.scala 90:30]
  assign _T_1594 = _T_1591[15:0]; // @[Shift.scala 90:48]
  assign _T_1595 = _T_1594 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_22 = {{16'd0}, _T_1595}; // @[Shift.scala 90:39]
  assign _T_1596 = _T_1593 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_1597 = _T_1592[4]; // @[Shift.scala 12:21]
  assign _T_1598 = _T_1591[32]; // @[Shift.scala 12:21]
  assign _T_1600 = _T_1598 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_1601 = {_T_1600,_T_1596}; // @[Cat.scala 29:58]
  assign _T_1602 = _T_1597 ? _T_1601 : _T_1591; // @[Shift.scala 91:22]
  assign _T_1603 = _T_1592[3:0]; // @[Shift.scala 92:77]
  assign _T_1604 = _T_1602[32:8]; // @[Shift.scala 90:30]
  assign _T_1605 = _T_1602[7:0]; // @[Shift.scala 90:48]
  assign _T_1606 = _T_1605 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_23 = {{24'd0}, _T_1606}; // @[Shift.scala 90:39]
  assign _T_1607 = _T_1604 | _GEN_23; // @[Shift.scala 90:39]
  assign _T_1608 = _T_1603[3]; // @[Shift.scala 12:21]
  assign _T_1609 = _T_1602[32]; // @[Shift.scala 12:21]
  assign _T_1611 = _T_1609 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_1612 = {_T_1611,_T_1607}; // @[Cat.scala 29:58]
  assign _T_1613 = _T_1608 ? _T_1612 : _T_1602; // @[Shift.scala 91:22]
  assign _T_1614 = _T_1603[2:0]; // @[Shift.scala 92:77]
  assign _T_1615 = _T_1613[32:4]; // @[Shift.scala 90:30]
  assign _T_1616 = _T_1613[3:0]; // @[Shift.scala 90:48]
  assign _T_1617 = _T_1616 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_24 = {{28'd0}, _T_1617}; // @[Shift.scala 90:39]
  assign _T_1618 = _T_1615 | _GEN_24; // @[Shift.scala 90:39]
  assign _T_1619 = _T_1614[2]; // @[Shift.scala 12:21]
  assign _T_1620 = _T_1613[32]; // @[Shift.scala 12:21]
  assign _T_1622 = _T_1620 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_1623 = {_T_1622,_T_1618}; // @[Cat.scala 29:58]
  assign _T_1624 = _T_1619 ? _T_1623 : _T_1613; // @[Shift.scala 91:22]
  assign _T_1625 = _T_1614[1:0]; // @[Shift.scala 92:77]
  assign _T_1626 = _T_1624[32:2]; // @[Shift.scala 90:30]
  assign _T_1627 = _T_1624[1:0]; // @[Shift.scala 90:48]
  assign _T_1628 = _T_1627 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_25 = {{30'd0}, _T_1628}; // @[Shift.scala 90:39]
  assign _T_1629 = _T_1626 | _GEN_25; // @[Shift.scala 90:39]
  assign _T_1630 = _T_1625[1]; // @[Shift.scala 12:21]
  assign _T_1631 = _T_1624[32]; // @[Shift.scala 12:21]
  assign _T_1633 = _T_1631 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_1634 = {_T_1633,_T_1629}; // @[Cat.scala 29:58]
  assign _T_1635 = _T_1630 ? _T_1634 : _T_1624; // @[Shift.scala 91:22]
  assign _T_1636 = _T_1625[0:0]; // @[Shift.scala 92:77]
  assign _T_1637 = _T_1635[32:1]; // @[Shift.scala 90:30]
  assign _T_1638 = _T_1635[0:0]; // @[Shift.scala 90:48]
  assign _GEN_26 = {{31'd0}, _T_1638}; // @[Shift.scala 90:39]
  assign _T_1640 = _T_1637 | _GEN_26; // @[Shift.scala 90:39]
  assign _T_1642 = _T_1635[32]; // @[Shift.scala 12:21]
  assign _T_1643 = {_T_1642,_T_1640}; // @[Cat.scala 29:58]
  assign _T_1644 = _T_1636 ? _T_1643 : _T_1635; // @[Shift.scala 91:22]
  assign _T_1647 = _T_1587 ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 71:12]
  assign _T_1648 = _T_1580 ? _T_1644 : _T_1647; // @[Shift.scala 39:10]
  assign _T_1649 = _T_1648[3]; // @[convert.scala 55:31]
  assign _T_1650 = _T_1648[2]; // @[convert.scala 56:31]
  assign _T_1651 = _T_1648[1]; // @[convert.scala 57:31]
  assign _T_1652 = _T_1648[0]; // @[convert.scala 58:31]
  assign _T_1653 = _T_1648[32:3]; // @[convert.scala 59:69]
  assign _T_1654 = _T_1653 != 30'h0; // @[convert.scala 59:81]
  assign _T_1655 = ~ _T_1654; // @[convert.scala 59:50]
  assign _T_1657 = _T_1653 == 30'h3fffffff; // @[convert.scala 60:81]
  assign _T_1658 = _T_1649 | _T_1651; // @[convert.scala 61:44]
  assign _T_1659 = _T_1658 | _T_1652; // @[convert.scala 61:52]
  assign _T_1660 = _T_1650 & _T_1659; // @[convert.scala 61:36]
  assign _T_1661 = ~ _T_1657; // @[convert.scala 62:63]
  assign _T_1662 = _T_1661 & _T_1660; // @[convert.scala 62:103]
  assign _T_1663 = _T_1655 | _T_1662; // @[convert.scala 62:60]
  assign _GEN_27 = {{29'd0}, _T_1663}; // @[convert.scala 63:56]
  assign _T_1666 = _T_1653 + _GEN_27; // @[convert.scala 63:56]
  assign _T_1667 = {sumSign,_T_1666}; // @[Cat.scala 29:58]
  assign io_F = _T_1675; // @[PositFMA.scala 174:15]
  assign io_outValid = _T_1671; // @[PositFMA.scala 173:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  outIsNaR_phase2 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  mulSig_phase2 = _RAND_1[52:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  addFrac_phase2 = _RAND_2[24:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mulScale_phase2 = _RAND_3[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addScale_phase2 = _RAND_4[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addSign_phase2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addZero_phase2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  inValid_phase2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1671 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_1675 = _RAND_9[30:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (io_inValid) begin
      outIsNaR_phase2 <= outIsNaR;
    end
    if (io_inValid) begin
      mulSig_phase2 <= mulSig;
    end
    if (io_inValid) begin
      addFrac_phase2 <= decC_fraction;
    end
    if (io_inValid) begin
      mulScale_phase2 <= mulScale;
    end
    if (io_inValid) begin
      addScale_phase2 <= decC_scale;
    end
    if (io_inValid) begin
      addSign_phase2 <= _T_619;
    end
    if (io_inValid) begin
      addZero_phase2 <= decC_isZero;
    end
    if (reset) begin
      inValid_phase2 <= 1'h0;
    end else begin
      inValid_phase2 <= io_inValid;
    end
    if (reset) begin
      _T_1671 <= 1'h0;
    end else begin
      _T_1671 <= inValid_phase2;
    end
    if (inValid_phase2) begin
      if (outIsNaR_phase2) begin
        _T_1675 <= 31'h40000000;
      end else begin
        if (decF_isZero) begin
          _T_1675 <= 31'h0;
        end else begin
          _T_1675 <= _T_1667;
        end
      end
    end
  end
endmodule
