module PositMultiplier28_3(
  input         clock,
  input         reset,
  input  [27:0] io_A,
  input  [27:0] io_B,
  output [27:0] io_M
);
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [25:0] _T_4; // @[convert.scala 19:24]
  wire [25:0] _T_5; // @[convert.scala 19:43]
  wire [25:0] _T_6; // @[convert.scala 19:39]
  wire [15:0] _T_7; // @[LZD.scala 43:32]
  wire [7:0] _T_8; // @[LZD.scala 43:32]
  wire [3:0] _T_9; // @[LZD.scala 43:32]
  wire [1:0] _T_10; // @[LZD.scala 43:32]
  wire  _T_11; // @[LZD.scala 39:14]
  wire  _T_12; // @[LZD.scala 39:21]
  wire  _T_13; // @[LZD.scala 39:30]
  wire  _T_14; // @[LZD.scala 39:27]
  wire  _T_15; // @[LZD.scala 39:25]
  wire [1:0] _T_16; // @[Cat.scala 29:58]
  wire [1:0] _T_17; // @[LZD.scala 44:32]
  wire  _T_18; // @[LZD.scala 39:14]
  wire  _T_19; // @[LZD.scala 39:21]
  wire  _T_20; // @[LZD.scala 39:30]
  wire  _T_21; // @[LZD.scala 39:27]
  wire  _T_22; // @[LZD.scala 39:25]
  wire [1:0] _T_23; // @[Cat.scala 29:58]
  wire  _T_24; // @[Shift.scala 12:21]
  wire  _T_25; // @[Shift.scala 12:21]
  wire  _T_26; // @[LZD.scala 49:16]
  wire  _T_27; // @[LZD.scala 49:27]
  wire  _T_28; // @[LZD.scala 49:25]
  wire  _T_29; // @[LZD.scala 49:47]
  wire  _T_30; // @[LZD.scala 49:59]
  wire  _T_31; // @[LZD.scala 49:35]
  wire [2:0] _T_33; // @[Cat.scala 29:58]
  wire [3:0] _T_34; // @[LZD.scala 44:32]
  wire [1:0] _T_35; // @[LZD.scala 43:32]
  wire  _T_36; // @[LZD.scala 39:14]
  wire  _T_37; // @[LZD.scala 39:21]
  wire  _T_38; // @[LZD.scala 39:30]
  wire  _T_39; // @[LZD.scala 39:27]
  wire  _T_40; // @[LZD.scala 39:25]
  wire [1:0] _T_41; // @[Cat.scala 29:58]
  wire [1:0] _T_42; // @[LZD.scala 44:32]
  wire  _T_43; // @[LZD.scala 39:14]
  wire  _T_44; // @[LZD.scala 39:21]
  wire  _T_45; // @[LZD.scala 39:30]
  wire  _T_46; // @[LZD.scala 39:27]
  wire  _T_47; // @[LZD.scala 39:25]
  wire [1:0] _T_48; // @[Cat.scala 29:58]
  wire  _T_49; // @[Shift.scala 12:21]
  wire  _T_50; // @[Shift.scala 12:21]
  wire  _T_51; // @[LZD.scala 49:16]
  wire  _T_52; // @[LZD.scala 49:27]
  wire  _T_53; // @[LZD.scala 49:25]
  wire  _T_54; // @[LZD.scala 49:47]
  wire  _T_55; // @[LZD.scala 49:59]
  wire  _T_56; // @[LZD.scala 49:35]
  wire [2:0] _T_58; // @[Cat.scala 29:58]
  wire  _T_59; // @[Shift.scala 12:21]
  wire  _T_60; // @[Shift.scala 12:21]
  wire  _T_61; // @[LZD.scala 49:16]
  wire  _T_62; // @[LZD.scala 49:27]
  wire  _T_63; // @[LZD.scala 49:25]
  wire [1:0] _T_64; // @[LZD.scala 49:47]
  wire [1:0] _T_65; // @[LZD.scala 49:59]
  wire [1:0] _T_66; // @[LZD.scala 49:35]
  wire [3:0] _T_68; // @[Cat.scala 29:58]
  wire [7:0] _T_69; // @[LZD.scala 44:32]
  wire [3:0] _T_70; // @[LZD.scala 43:32]
  wire [1:0] _T_71; // @[LZD.scala 43:32]
  wire  _T_72; // @[LZD.scala 39:14]
  wire  _T_73; // @[LZD.scala 39:21]
  wire  _T_74; // @[LZD.scala 39:30]
  wire  _T_75; // @[LZD.scala 39:27]
  wire  _T_76; // @[LZD.scala 39:25]
  wire [1:0] _T_77; // @[Cat.scala 29:58]
  wire [1:0] _T_78; // @[LZD.scala 44:32]
  wire  _T_79; // @[LZD.scala 39:14]
  wire  _T_80; // @[LZD.scala 39:21]
  wire  _T_81; // @[LZD.scala 39:30]
  wire  _T_82; // @[LZD.scala 39:27]
  wire  _T_83; // @[LZD.scala 39:25]
  wire [1:0] _T_84; // @[Cat.scala 29:58]
  wire  _T_85; // @[Shift.scala 12:21]
  wire  _T_86; // @[Shift.scala 12:21]
  wire  _T_87; // @[LZD.scala 49:16]
  wire  _T_88; // @[LZD.scala 49:27]
  wire  _T_89; // @[LZD.scala 49:25]
  wire  _T_90; // @[LZD.scala 49:47]
  wire  _T_91; // @[LZD.scala 49:59]
  wire  _T_92; // @[LZD.scala 49:35]
  wire [2:0] _T_94; // @[Cat.scala 29:58]
  wire [3:0] _T_95; // @[LZD.scala 44:32]
  wire [1:0] _T_96; // @[LZD.scala 43:32]
  wire  _T_97; // @[LZD.scala 39:14]
  wire  _T_98; // @[LZD.scala 39:21]
  wire  _T_99; // @[LZD.scala 39:30]
  wire  _T_100; // @[LZD.scala 39:27]
  wire  _T_101; // @[LZD.scala 39:25]
  wire [1:0] _T_102; // @[Cat.scala 29:58]
  wire [1:0] _T_103; // @[LZD.scala 44:32]
  wire  _T_104; // @[LZD.scala 39:14]
  wire  _T_105; // @[LZD.scala 39:21]
  wire  _T_106; // @[LZD.scala 39:30]
  wire  _T_107; // @[LZD.scala 39:27]
  wire  _T_108; // @[LZD.scala 39:25]
  wire [1:0] _T_109; // @[Cat.scala 29:58]
  wire  _T_110; // @[Shift.scala 12:21]
  wire  _T_111; // @[Shift.scala 12:21]
  wire  _T_112; // @[LZD.scala 49:16]
  wire  _T_113; // @[LZD.scala 49:27]
  wire  _T_114; // @[LZD.scala 49:25]
  wire  _T_115; // @[LZD.scala 49:47]
  wire  _T_116; // @[LZD.scala 49:59]
  wire  _T_117; // @[LZD.scala 49:35]
  wire [2:0] _T_119; // @[Cat.scala 29:58]
  wire  _T_120; // @[Shift.scala 12:21]
  wire  _T_121; // @[Shift.scala 12:21]
  wire  _T_122; // @[LZD.scala 49:16]
  wire  _T_123; // @[LZD.scala 49:27]
  wire  _T_124; // @[LZD.scala 49:25]
  wire [1:0] _T_125; // @[LZD.scala 49:47]
  wire [1:0] _T_126; // @[LZD.scala 49:59]
  wire [1:0] _T_127; // @[LZD.scala 49:35]
  wire [3:0] _T_129; // @[Cat.scala 29:58]
  wire  _T_130; // @[Shift.scala 12:21]
  wire  _T_131; // @[Shift.scala 12:21]
  wire  _T_132; // @[LZD.scala 49:16]
  wire  _T_133; // @[LZD.scala 49:27]
  wire  _T_134; // @[LZD.scala 49:25]
  wire [2:0] _T_135; // @[LZD.scala 49:47]
  wire [2:0] _T_136; // @[LZD.scala 49:59]
  wire [2:0] _T_137; // @[LZD.scala 49:35]
  wire [4:0] _T_139; // @[Cat.scala 29:58]
  wire [9:0] _T_140; // @[LZD.scala 44:32]
  wire [7:0] _T_141; // @[LZD.scala 43:32]
  wire [3:0] _T_142; // @[LZD.scala 43:32]
  wire [1:0] _T_143; // @[LZD.scala 43:32]
  wire  _T_144; // @[LZD.scala 39:14]
  wire  _T_145; // @[LZD.scala 39:21]
  wire  _T_146; // @[LZD.scala 39:30]
  wire  _T_147; // @[LZD.scala 39:27]
  wire  _T_148; // @[LZD.scala 39:25]
  wire [1:0] _T_149; // @[Cat.scala 29:58]
  wire [1:0] _T_150; // @[LZD.scala 44:32]
  wire  _T_151; // @[LZD.scala 39:14]
  wire  _T_152; // @[LZD.scala 39:21]
  wire  _T_153; // @[LZD.scala 39:30]
  wire  _T_154; // @[LZD.scala 39:27]
  wire  _T_155; // @[LZD.scala 39:25]
  wire [1:0] _T_156; // @[Cat.scala 29:58]
  wire  _T_157; // @[Shift.scala 12:21]
  wire  _T_158; // @[Shift.scala 12:21]
  wire  _T_159; // @[LZD.scala 49:16]
  wire  _T_160; // @[LZD.scala 49:27]
  wire  _T_161; // @[LZD.scala 49:25]
  wire  _T_162; // @[LZD.scala 49:47]
  wire  _T_163; // @[LZD.scala 49:59]
  wire  _T_164; // @[LZD.scala 49:35]
  wire [2:0] _T_166; // @[Cat.scala 29:58]
  wire [3:0] _T_167; // @[LZD.scala 44:32]
  wire [1:0] _T_168; // @[LZD.scala 43:32]
  wire  _T_169; // @[LZD.scala 39:14]
  wire  _T_170; // @[LZD.scala 39:21]
  wire  _T_171; // @[LZD.scala 39:30]
  wire  _T_172; // @[LZD.scala 39:27]
  wire  _T_173; // @[LZD.scala 39:25]
  wire [1:0] _T_174; // @[Cat.scala 29:58]
  wire [1:0] _T_175; // @[LZD.scala 44:32]
  wire  _T_176; // @[LZD.scala 39:14]
  wire  _T_177; // @[LZD.scala 39:21]
  wire  _T_178; // @[LZD.scala 39:30]
  wire  _T_179; // @[LZD.scala 39:27]
  wire  _T_180; // @[LZD.scala 39:25]
  wire [1:0] _T_181; // @[Cat.scala 29:58]
  wire  _T_182; // @[Shift.scala 12:21]
  wire  _T_183; // @[Shift.scala 12:21]
  wire  _T_184; // @[LZD.scala 49:16]
  wire  _T_185; // @[LZD.scala 49:27]
  wire  _T_186; // @[LZD.scala 49:25]
  wire  _T_187; // @[LZD.scala 49:47]
  wire  _T_188; // @[LZD.scala 49:59]
  wire  _T_189; // @[LZD.scala 49:35]
  wire [2:0] _T_191; // @[Cat.scala 29:58]
  wire  _T_192; // @[Shift.scala 12:21]
  wire  _T_193; // @[Shift.scala 12:21]
  wire  _T_194; // @[LZD.scala 49:16]
  wire  _T_195; // @[LZD.scala 49:27]
  wire  _T_196; // @[LZD.scala 49:25]
  wire [1:0] _T_197; // @[LZD.scala 49:47]
  wire [1:0] _T_198; // @[LZD.scala 49:59]
  wire [1:0] _T_199; // @[LZD.scala 49:35]
  wire [3:0] _T_201; // @[Cat.scala 29:58]
  wire [1:0] _T_202; // @[LZD.scala 44:32]
  wire  _T_203; // @[LZD.scala 39:14]
  wire  _T_204; // @[LZD.scala 39:21]
  wire  _T_205; // @[LZD.scala 39:30]
  wire  _T_206; // @[LZD.scala 39:27]
  wire  _T_207; // @[LZD.scala 39:25]
  wire  _T_209; // @[Shift.scala 12:21]
  wire [2:0] _T_211; // @[Cat.scala 29:58]
  wire [2:0] _T_212; // @[LZD.scala 55:32]
  wire [2:0] _T_213; // @[LZD.scala 55:20]
  wire [3:0] _T_214; // @[Cat.scala 29:58]
  wire  _T_215; // @[Shift.scala 12:21]
  wire [3:0] _T_217; // @[LZD.scala 55:32]
  wire [3:0] _T_218; // @[LZD.scala 55:20]
  wire [4:0] _T_219; // @[Cat.scala 29:58]
  wire [4:0] _T_220; // @[convert.scala 21:22]
  wire [24:0] _T_221; // @[convert.scala 22:36]
  wire  _T_222; // @[Shift.scala 16:24]
  wire  _T_224; // @[Shift.scala 12:21]
  wire [8:0] _T_225; // @[Shift.scala 64:52]
  wire [24:0] _T_227; // @[Cat.scala 29:58]
  wire [24:0] _T_228; // @[Shift.scala 64:27]
  wire [3:0] _T_229; // @[Shift.scala 66:70]
  wire  _T_230; // @[Shift.scala 12:21]
  wire [16:0] _T_231; // @[Shift.scala 64:52]
  wire [24:0] _T_233; // @[Cat.scala 29:58]
  wire [24:0] _T_234; // @[Shift.scala 64:27]
  wire [2:0] _T_235; // @[Shift.scala 66:70]
  wire  _T_236; // @[Shift.scala 12:21]
  wire [20:0] _T_237; // @[Shift.scala 64:52]
  wire [24:0] _T_239; // @[Cat.scala 29:58]
  wire [24:0] _T_240; // @[Shift.scala 64:27]
  wire [1:0] _T_241; // @[Shift.scala 66:70]
  wire  _T_242; // @[Shift.scala 12:21]
  wire [22:0] _T_243; // @[Shift.scala 64:52]
  wire [24:0] _T_245; // @[Cat.scala 29:58]
  wire [24:0] _T_246; // @[Shift.scala 64:27]
  wire  _T_247; // @[Shift.scala 66:70]
  wire [23:0] _T_249; // @[Shift.scala 64:52]
  wire [24:0] _T_250; // @[Cat.scala 29:58]
  wire [24:0] _T_251; // @[Shift.scala 64:27]
  wire [24:0] _T_252; // @[Shift.scala 16:10]
  wire [2:0] _T_253; // @[convert.scala 23:34]
  wire [21:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_255; // @[convert.scala 25:26]
  wire [4:0] _T_257; // @[convert.scala 25:42]
  wire [2:0] _T_260; // @[convert.scala 26:67]
  wire [2:0] _T_261; // @[convert.scala 26:51]
  wire [8:0] _T_262; // @[Cat.scala 29:58]
  wire [26:0] _T_264; // @[convert.scala 29:56]
  wire  _T_265; // @[convert.scala 29:60]
  wire  _T_266; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_269; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [8:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_278; // @[convert.scala 18:24]
  wire  _T_279; // @[convert.scala 18:40]
  wire  _T_280; // @[convert.scala 18:36]
  wire [25:0] _T_281; // @[convert.scala 19:24]
  wire [25:0] _T_282; // @[convert.scala 19:43]
  wire [25:0] _T_283; // @[convert.scala 19:39]
  wire [15:0] _T_284; // @[LZD.scala 43:32]
  wire [7:0] _T_285; // @[LZD.scala 43:32]
  wire [3:0] _T_286; // @[LZD.scala 43:32]
  wire [1:0] _T_287; // @[LZD.scala 43:32]
  wire  _T_288; // @[LZD.scala 39:14]
  wire  _T_289; // @[LZD.scala 39:21]
  wire  _T_290; // @[LZD.scala 39:30]
  wire  _T_291; // @[LZD.scala 39:27]
  wire  _T_292; // @[LZD.scala 39:25]
  wire [1:0] _T_293; // @[Cat.scala 29:58]
  wire [1:0] _T_294; // @[LZD.scala 44:32]
  wire  _T_295; // @[LZD.scala 39:14]
  wire  _T_296; // @[LZD.scala 39:21]
  wire  _T_297; // @[LZD.scala 39:30]
  wire  _T_298; // @[LZD.scala 39:27]
  wire  _T_299; // @[LZD.scala 39:25]
  wire [1:0] _T_300; // @[Cat.scala 29:58]
  wire  _T_301; // @[Shift.scala 12:21]
  wire  _T_302; // @[Shift.scala 12:21]
  wire  _T_303; // @[LZD.scala 49:16]
  wire  _T_304; // @[LZD.scala 49:27]
  wire  _T_305; // @[LZD.scala 49:25]
  wire  _T_306; // @[LZD.scala 49:47]
  wire  _T_307; // @[LZD.scala 49:59]
  wire  _T_308; // @[LZD.scala 49:35]
  wire [2:0] _T_310; // @[Cat.scala 29:58]
  wire [3:0] _T_311; // @[LZD.scala 44:32]
  wire [1:0] _T_312; // @[LZD.scala 43:32]
  wire  _T_313; // @[LZD.scala 39:14]
  wire  _T_314; // @[LZD.scala 39:21]
  wire  _T_315; // @[LZD.scala 39:30]
  wire  _T_316; // @[LZD.scala 39:27]
  wire  _T_317; // @[LZD.scala 39:25]
  wire [1:0] _T_318; // @[Cat.scala 29:58]
  wire [1:0] _T_319; // @[LZD.scala 44:32]
  wire  _T_320; // @[LZD.scala 39:14]
  wire  _T_321; // @[LZD.scala 39:21]
  wire  _T_322; // @[LZD.scala 39:30]
  wire  _T_323; // @[LZD.scala 39:27]
  wire  _T_324; // @[LZD.scala 39:25]
  wire [1:0] _T_325; // @[Cat.scala 29:58]
  wire  _T_326; // @[Shift.scala 12:21]
  wire  _T_327; // @[Shift.scala 12:21]
  wire  _T_328; // @[LZD.scala 49:16]
  wire  _T_329; // @[LZD.scala 49:27]
  wire  _T_330; // @[LZD.scala 49:25]
  wire  _T_331; // @[LZD.scala 49:47]
  wire  _T_332; // @[LZD.scala 49:59]
  wire  _T_333; // @[LZD.scala 49:35]
  wire [2:0] _T_335; // @[Cat.scala 29:58]
  wire  _T_336; // @[Shift.scala 12:21]
  wire  _T_337; // @[Shift.scala 12:21]
  wire  _T_338; // @[LZD.scala 49:16]
  wire  _T_339; // @[LZD.scala 49:27]
  wire  _T_340; // @[LZD.scala 49:25]
  wire [1:0] _T_341; // @[LZD.scala 49:47]
  wire [1:0] _T_342; // @[LZD.scala 49:59]
  wire [1:0] _T_343; // @[LZD.scala 49:35]
  wire [3:0] _T_345; // @[Cat.scala 29:58]
  wire [7:0] _T_346; // @[LZD.scala 44:32]
  wire [3:0] _T_347; // @[LZD.scala 43:32]
  wire [1:0] _T_348; // @[LZD.scala 43:32]
  wire  _T_349; // @[LZD.scala 39:14]
  wire  _T_350; // @[LZD.scala 39:21]
  wire  _T_351; // @[LZD.scala 39:30]
  wire  _T_352; // @[LZD.scala 39:27]
  wire  _T_353; // @[LZD.scala 39:25]
  wire [1:0] _T_354; // @[Cat.scala 29:58]
  wire [1:0] _T_355; // @[LZD.scala 44:32]
  wire  _T_356; // @[LZD.scala 39:14]
  wire  _T_357; // @[LZD.scala 39:21]
  wire  _T_358; // @[LZD.scala 39:30]
  wire  _T_359; // @[LZD.scala 39:27]
  wire  _T_360; // @[LZD.scala 39:25]
  wire [1:0] _T_361; // @[Cat.scala 29:58]
  wire  _T_362; // @[Shift.scala 12:21]
  wire  _T_363; // @[Shift.scala 12:21]
  wire  _T_364; // @[LZD.scala 49:16]
  wire  _T_365; // @[LZD.scala 49:27]
  wire  _T_366; // @[LZD.scala 49:25]
  wire  _T_367; // @[LZD.scala 49:47]
  wire  _T_368; // @[LZD.scala 49:59]
  wire  _T_369; // @[LZD.scala 49:35]
  wire [2:0] _T_371; // @[Cat.scala 29:58]
  wire [3:0] _T_372; // @[LZD.scala 44:32]
  wire [1:0] _T_373; // @[LZD.scala 43:32]
  wire  _T_374; // @[LZD.scala 39:14]
  wire  _T_375; // @[LZD.scala 39:21]
  wire  _T_376; // @[LZD.scala 39:30]
  wire  _T_377; // @[LZD.scala 39:27]
  wire  _T_378; // @[LZD.scala 39:25]
  wire [1:0] _T_379; // @[Cat.scala 29:58]
  wire [1:0] _T_380; // @[LZD.scala 44:32]
  wire  _T_381; // @[LZD.scala 39:14]
  wire  _T_382; // @[LZD.scala 39:21]
  wire  _T_383; // @[LZD.scala 39:30]
  wire  _T_384; // @[LZD.scala 39:27]
  wire  _T_385; // @[LZD.scala 39:25]
  wire [1:0] _T_386; // @[Cat.scala 29:58]
  wire  _T_387; // @[Shift.scala 12:21]
  wire  _T_388; // @[Shift.scala 12:21]
  wire  _T_389; // @[LZD.scala 49:16]
  wire  _T_390; // @[LZD.scala 49:27]
  wire  _T_391; // @[LZD.scala 49:25]
  wire  _T_392; // @[LZD.scala 49:47]
  wire  _T_393; // @[LZD.scala 49:59]
  wire  _T_394; // @[LZD.scala 49:35]
  wire [2:0] _T_396; // @[Cat.scala 29:58]
  wire  _T_397; // @[Shift.scala 12:21]
  wire  _T_398; // @[Shift.scala 12:21]
  wire  _T_399; // @[LZD.scala 49:16]
  wire  _T_400; // @[LZD.scala 49:27]
  wire  _T_401; // @[LZD.scala 49:25]
  wire [1:0] _T_402; // @[LZD.scala 49:47]
  wire [1:0] _T_403; // @[LZD.scala 49:59]
  wire [1:0] _T_404; // @[LZD.scala 49:35]
  wire [3:0] _T_406; // @[Cat.scala 29:58]
  wire  _T_407; // @[Shift.scala 12:21]
  wire  _T_408; // @[Shift.scala 12:21]
  wire  _T_409; // @[LZD.scala 49:16]
  wire  _T_410; // @[LZD.scala 49:27]
  wire  _T_411; // @[LZD.scala 49:25]
  wire [2:0] _T_412; // @[LZD.scala 49:47]
  wire [2:0] _T_413; // @[LZD.scala 49:59]
  wire [2:0] _T_414; // @[LZD.scala 49:35]
  wire [4:0] _T_416; // @[Cat.scala 29:58]
  wire [9:0] _T_417; // @[LZD.scala 44:32]
  wire [7:0] _T_418; // @[LZD.scala 43:32]
  wire [3:0] _T_419; // @[LZD.scala 43:32]
  wire [1:0] _T_420; // @[LZD.scala 43:32]
  wire  _T_421; // @[LZD.scala 39:14]
  wire  _T_422; // @[LZD.scala 39:21]
  wire  _T_423; // @[LZD.scala 39:30]
  wire  _T_424; // @[LZD.scala 39:27]
  wire  _T_425; // @[LZD.scala 39:25]
  wire [1:0] _T_426; // @[Cat.scala 29:58]
  wire [1:0] _T_427; // @[LZD.scala 44:32]
  wire  _T_428; // @[LZD.scala 39:14]
  wire  _T_429; // @[LZD.scala 39:21]
  wire  _T_430; // @[LZD.scala 39:30]
  wire  _T_431; // @[LZD.scala 39:27]
  wire  _T_432; // @[LZD.scala 39:25]
  wire [1:0] _T_433; // @[Cat.scala 29:58]
  wire  _T_434; // @[Shift.scala 12:21]
  wire  _T_435; // @[Shift.scala 12:21]
  wire  _T_436; // @[LZD.scala 49:16]
  wire  _T_437; // @[LZD.scala 49:27]
  wire  _T_438; // @[LZD.scala 49:25]
  wire  _T_439; // @[LZD.scala 49:47]
  wire  _T_440; // @[LZD.scala 49:59]
  wire  _T_441; // @[LZD.scala 49:35]
  wire [2:0] _T_443; // @[Cat.scala 29:58]
  wire [3:0] _T_444; // @[LZD.scala 44:32]
  wire [1:0] _T_445; // @[LZD.scala 43:32]
  wire  _T_446; // @[LZD.scala 39:14]
  wire  _T_447; // @[LZD.scala 39:21]
  wire  _T_448; // @[LZD.scala 39:30]
  wire  _T_449; // @[LZD.scala 39:27]
  wire  _T_450; // @[LZD.scala 39:25]
  wire [1:0] _T_451; // @[Cat.scala 29:58]
  wire [1:0] _T_452; // @[LZD.scala 44:32]
  wire  _T_453; // @[LZD.scala 39:14]
  wire  _T_454; // @[LZD.scala 39:21]
  wire  _T_455; // @[LZD.scala 39:30]
  wire  _T_456; // @[LZD.scala 39:27]
  wire  _T_457; // @[LZD.scala 39:25]
  wire [1:0] _T_458; // @[Cat.scala 29:58]
  wire  _T_459; // @[Shift.scala 12:21]
  wire  _T_460; // @[Shift.scala 12:21]
  wire  _T_461; // @[LZD.scala 49:16]
  wire  _T_462; // @[LZD.scala 49:27]
  wire  _T_463; // @[LZD.scala 49:25]
  wire  _T_464; // @[LZD.scala 49:47]
  wire  _T_465; // @[LZD.scala 49:59]
  wire  _T_466; // @[LZD.scala 49:35]
  wire [2:0] _T_468; // @[Cat.scala 29:58]
  wire  _T_469; // @[Shift.scala 12:21]
  wire  _T_470; // @[Shift.scala 12:21]
  wire  _T_471; // @[LZD.scala 49:16]
  wire  _T_472; // @[LZD.scala 49:27]
  wire  _T_473; // @[LZD.scala 49:25]
  wire [1:0] _T_474; // @[LZD.scala 49:47]
  wire [1:0] _T_475; // @[LZD.scala 49:59]
  wire [1:0] _T_476; // @[LZD.scala 49:35]
  wire [3:0] _T_478; // @[Cat.scala 29:58]
  wire [1:0] _T_479; // @[LZD.scala 44:32]
  wire  _T_480; // @[LZD.scala 39:14]
  wire  _T_481; // @[LZD.scala 39:21]
  wire  _T_482; // @[LZD.scala 39:30]
  wire  _T_483; // @[LZD.scala 39:27]
  wire  _T_484; // @[LZD.scala 39:25]
  wire  _T_486; // @[Shift.scala 12:21]
  wire [2:0] _T_488; // @[Cat.scala 29:58]
  wire [2:0] _T_489; // @[LZD.scala 55:32]
  wire [2:0] _T_490; // @[LZD.scala 55:20]
  wire [3:0] _T_491; // @[Cat.scala 29:58]
  wire  _T_492; // @[Shift.scala 12:21]
  wire [3:0] _T_494; // @[LZD.scala 55:32]
  wire [3:0] _T_495; // @[LZD.scala 55:20]
  wire [4:0] _T_496; // @[Cat.scala 29:58]
  wire [4:0] _T_497; // @[convert.scala 21:22]
  wire [24:0] _T_498; // @[convert.scala 22:36]
  wire  _T_499; // @[Shift.scala 16:24]
  wire  _T_501; // @[Shift.scala 12:21]
  wire [8:0] _T_502; // @[Shift.scala 64:52]
  wire [24:0] _T_504; // @[Cat.scala 29:58]
  wire [24:0] _T_505; // @[Shift.scala 64:27]
  wire [3:0] _T_506; // @[Shift.scala 66:70]
  wire  _T_507; // @[Shift.scala 12:21]
  wire [16:0] _T_508; // @[Shift.scala 64:52]
  wire [24:0] _T_510; // @[Cat.scala 29:58]
  wire [24:0] _T_511; // @[Shift.scala 64:27]
  wire [2:0] _T_512; // @[Shift.scala 66:70]
  wire  _T_513; // @[Shift.scala 12:21]
  wire [20:0] _T_514; // @[Shift.scala 64:52]
  wire [24:0] _T_516; // @[Cat.scala 29:58]
  wire [24:0] _T_517; // @[Shift.scala 64:27]
  wire [1:0] _T_518; // @[Shift.scala 66:70]
  wire  _T_519; // @[Shift.scala 12:21]
  wire [22:0] _T_520; // @[Shift.scala 64:52]
  wire [24:0] _T_522; // @[Cat.scala 29:58]
  wire [24:0] _T_523; // @[Shift.scala 64:27]
  wire  _T_524; // @[Shift.scala 66:70]
  wire [23:0] _T_526; // @[Shift.scala 64:52]
  wire [24:0] _T_527; // @[Cat.scala 29:58]
  wire [24:0] _T_528; // @[Shift.scala 64:27]
  wire [24:0] _T_529; // @[Shift.scala 16:10]
  wire [2:0] _T_530; // @[convert.scala 23:34]
  wire [21:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_532; // @[convert.scala 25:26]
  wire [4:0] _T_534; // @[convert.scala 25:42]
  wire [2:0] _T_537; // @[convert.scala 26:67]
  wire [2:0] _T_538; // @[convert.scala 26:51]
  wire [8:0] _T_539; // @[Cat.scala 29:58]
  wire [26:0] _T_541; // @[convert.scala 29:56]
  wire  _T_542; // @[convert.scala 29:60]
  wire  _T_543; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_546; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [8:0] decB_scale; // @[convert.scala 32:24]
  wire  _T_554; // @[PositMultiplier.scala 43:34]
  wire [23:0] _T_556; // @[Cat.scala 29:58]
  wire [23:0] sigA; // @[PositMultiplier.scala 43:61]
  wire  _T_557; // @[PositMultiplier.scala 44:34]
  wire [23:0] _T_559; // @[Cat.scala 29:58]
  wire [23:0] sigB; // @[PositMultiplier.scala 44:61]
  wire [47:0] _T_560; // @[PositMultiplier.scala 45:25]
  wire [47:0] sigP; // @[PositMultiplier.scala 45:33]
  wire [1:0] head2; // @[PositMultiplier.scala 46:28]
  wire  _T_561; // @[PositMultiplier.scala 47:31]
  wire  _T_562; // @[PositMultiplier.scala 47:25]
  wire  _T_563; // @[PositMultiplier.scala 47:42]
  wire  addTwo; // @[PositMultiplier.scala 47:35]
  wire  _T_564; // @[PositMultiplier.scala 49:23]
  wire  _T_565; // @[PositMultiplier.scala 49:49]
  wire  addOne; // @[PositMultiplier.scala 49:43]
  wire [1:0] _T_566; // @[Cat.scala 29:58]
  wire [2:0] expBias; // @[PositMultiplier.scala 50:39]
  wire [44:0] _T_567; // @[PositMultiplier.scala 53:81]
  wire [43:0] _T_568; // @[PositMultiplier.scala 54:81]
  wire [44:0] _T_569; // @[PositMultiplier.scala 54:104]
  wire [44:0] frac; // @[PositMultiplier.scala 51:22]
  wire [9:0] _T_570; // @[PositMultiplier.scala 56:30]
  wire [9:0] _GEN_0; // @[PositMultiplier.scala 56:44]
  wire [9:0] _T_572; // @[PositMultiplier.scala 56:44]
  wire [9:0] mulScale; // @[PositMultiplier.scala 56:44]
  wire  underflow; // @[PositMultiplier.scala 57:28]
  wire  overflow; // @[PositMultiplier.scala 58:28]
  wire  decM_sign; // @[PositMultiplier.scala 62:29]
  wire [9:0] _T_575; // @[Mux.scala 87:16]
  wire [9:0] _T_576; // @[Mux.scala 87:16]
  wire [21:0] decM_fraction; // @[PositMultiplier.scala 70:29]
  wire  decM_isNaR; // @[PositMultiplier.scala 71:31]
  wire  decM_isZero; // @[PositMultiplier.scala 72:32]
  wire [22:0] grsTmp; // @[PositMultiplier.scala 75:30]
  wire [1:0] _T_580; // @[PositMultiplier.scala 78:32]
  wire [20:0] _T_581; // @[PositMultiplier.scala 78:48]
  wire  _T_582; // @[PositMultiplier.scala 78:52]
  wire [8:0] _GEN_1; // @[PositMultiplier.scala 60:23 PositMultiplier.scala 63:17]
  wire [8:0] decM_scale; // @[PositMultiplier.scala 60:23 PositMultiplier.scala 63:17]
  wire [2:0] _T_585; // @[convert.scala 46:61]
  wire [2:0] _T_586; // @[convert.scala 46:52]
  wire [2:0] _T_588; // @[convert.scala 46:42]
  wire [5:0] _T_589; // @[convert.scala 48:34]
  wire  _T_590; // @[convert.scala 49:36]
  wire [5:0] _T_592; // @[convert.scala 50:36]
  wire [5:0] _T_593; // @[convert.scala 50:36]
  wire [5:0] _T_594; // @[convert.scala 50:28]
  wire  _T_595; // @[convert.scala 51:31]
  wire  _T_596; // @[convert.scala 52:43]
  wire [29:0] _T_600; // @[Cat.scala 29:58]
  wire [5:0] _T_601; // @[Shift.scala 39:17]
  wire  _T_602; // @[Shift.scala 39:24]
  wire [4:0] _T_603; // @[Shift.scala 40:44]
  wire [13:0] _T_604; // @[Shift.scala 90:30]
  wire [15:0] _T_605; // @[Shift.scala 90:48]
  wire  _T_606; // @[Shift.scala 90:57]
  wire [13:0] _GEN_2; // @[Shift.scala 90:39]
  wire [13:0] _T_607; // @[Shift.scala 90:39]
  wire  _T_608; // @[Shift.scala 12:21]
  wire  _T_609; // @[Shift.scala 12:21]
  wire [15:0] _T_611; // @[Bitwise.scala 71:12]
  wire [29:0] _T_612; // @[Cat.scala 29:58]
  wire [29:0] _T_613; // @[Shift.scala 91:22]
  wire [3:0] _T_614; // @[Shift.scala 92:77]
  wire [21:0] _T_615; // @[Shift.scala 90:30]
  wire [7:0] _T_616; // @[Shift.scala 90:48]
  wire  _T_617; // @[Shift.scala 90:57]
  wire [21:0] _GEN_3; // @[Shift.scala 90:39]
  wire [21:0] _T_618; // @[Shift.scala 90:39]
  wire  _T_619; // @[Shift.scala 12:21]
  wire  _T_620; // @[Shift.scala 12:21]
  wire [7:0] _T_622; // @[Bitwise.scala 71:12]
  wire [29:0] _T_623; // @[Cat.scala 29:58]
  wire [29:0] _T_624; // @[Shift.scala 91:22]
  wire [2:0] _T_625; // @[Shift.scala 92:77]
  wire [25:0] _T_626; // @[Shift.scala 90:30]
  wire [3:0] _T_627; // @[Shift.scala 90:48]
  wire  _T_628; // @[Shift.scala 90:57]
  wire [25:0] _GEN_4; // @[Shift.scala 90:39]
  wire [25:0] _T_629; // @[Shift.scala 90:39]
  wire  _T_630; // @[Shift.scala 12:21]
  wire  _T_631; // @[Shift.scala 12:21]
  wire [3:0] _T_633; // @[Bitwise.scala 71:12]
  wire [29:0] _T_634; // @[Cat.scala 29:58]
  wire [29:0] _T_635; // @[Shift.scala 91:22]
  wire [1:0] _T_636; // @[Shift.scala 92:77]
  wire [27:0] _T_637; // @[Shift.scala 90:30]
  wire [1:0] _T_638; // @[Shift.scala 90:48]
  wire  _T_639; // @[Shift.scala 90:57]
  wire [27:0] _GEN_5; // @[Shift.scala 90:39]
  wire [27:0] _T_640; // @[Shift.scala 90:39]
  wire  _T_641; // @[Shift.scala 12:21]
  wire  _T_642; // @[Shift.scala 12:21]
  wire [1:0] _T_644; // @[Bitwise.scala 71:12]
  wire [29:0] _T_645; // @[Cat.scala 29:58]
  wire [29:0] _T_646; // @[Shift.scala 91:22]
  wire  _T_647; // @[Shift.scala 92:77]
  wire [28:0] _T_648; // @[Shift.scala 90:30]
  wire  _T_649; // @[Shift.scala 90:48]
  wire [28:0] _GEN_6; // @[Shift.scala 90:39]
  wire [28:0] _T_651; // @[Shift.scala 90:39]
  wire  _T_653; // @[Shift.scala 12:21]
  wire [29:0] _T_654; // @[Cat.scala 29:58]
  wire [29:0] _T_655; // @[Shift.scala 91:22]
  wire [29:0] _T_658; // @[Bitwise.scala 71:12]
  wire [29:0] _T_659; // @[Shift.scala 39:10]
  wire  _T_660; // @[convert.scala 55:31]
  wire  _T_661; // @[convert.scala 56:31]
  wire  _T_662; // @[convert.scala 57:31]
  wire  _T_663; // @[convert.scala 58:31]
  wire [26:0] _T_664; // @[convert.scala 59:69]
  wire  _T_665; // @[convert.scala 59:81]
  wire  _T_666; // @[convert.scala 59:50]
  wire  _T_668; // @[convert.scala 60:81]
  wire  _T_669; // @[convert.scala 61:44]
  wire  _T_670; // @[convert.scala 61:52]
  wire  _T_671; // @[convert.scala 61:36]
  wire  _T_672; // @[convert.scala 62:63]
  wire  _T_673; // @[convert.scala 62:103]
  wire  _T_674; // @[convert.scala 62:60]
  wire [26:0] _GEN_7; // @[convert.scala 63:56]
  wire [26:0] _T_677; // @[convert.scala 63:56]
  wire [27:0] _T_678; // @[Cat.scala 29:58]
  wire [27:0] _T_680; // @[Mux.scala 87:16]
  assign _T_1 = io_A[27]; // @[convert.scala 18:24]
  assign _T_2 = io_A[26]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[26:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[25:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[25:10]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[15:8]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8[7:4]; // @[LZD.scala 43:32]
  assign _T_10 = _T_9[3:2]; // @[LZD.scala 43:32]
  assign _T_11 = _T_10 != 2'h0; // @[LZD.scala 39:14]
  assign _T_12 = _T_10[1]; // @[LZD.scala 39:21]
  assign _T_13 = _T_10[0]; // @[LZD.scala 39:30]
  assign _T_14 = ~ _T_13; // @[LZD.scala 39:27]
  assign _T_15 = _T_12 | _T_14; // @[LZD.scala 39:25]
  assign _T_16 = {_T_11,_T_15}; // @[Cat.scala 29:58]
  assign _T_17 = _T_9[1:0]; // @[LZD.scala 44:32]
  assign _T_18 = _T_17 != 2'h0; // @[LZD.scala 39:14]
  assign _T_19 = _T_17[1]; // @[LZD.scala 39:21]
  assign _T_20 = _T_17[0]; // @[LZD.scala 39:30]
  assign _T_21 = ~ _T_20; // @[LZD.scala 39:27]
  assign _T_22 = _T_19 | _T_21; // @[LZD.scala 39:25]
  assign _T_23 = {_T_18,_T_22}; // @[Cat.scala 29:58]
  assign _T_24 = _T_16[1]; // @[Shift.scala 12:21]
  assign _T_25 = _T_23[1]; // @[Shift.scala 12:21]
  assign _T_26 = _T_24 | _T_25; // @[LZD.scala 49:16]
  assign _T_27 = ~ _T_25; // @[LZD.scala 49:27]
  assign _T_28 = _T_24 | _T_27; // @[LZD.scala 49:25]
  assign _T_29 = _T_16[0:0]; // @[LZD.scala 49:47]
  assign _T_30 = _T_23[0:0]; // @[LZD.scala 49:59]
  assign _T_31 = _T_24 ? _T_29 : _T_30; // @[LZD.scala 49:35]
  assign _T_33 = {_T_26,_T_28,_T_31}; // @[Cat.scala 29:58]
  assign _T_34 = _T_8[3:0]; // @[LZD.scala 44:32]
  assign _T_35 = _T_34[3:2]; // @[LZD.scala 43:32]
  assign _T_36 = _T_35 != 2'h0; // @[LZD.scala 39:14]
  assign _T_37 = _T_35[1]; // @[LZD.scala 39:21]
  assign _T_38 = _T_35[0]; // @[LZD.scala 39:30]
  assign _T_39 = ~ _T_38; // @[LZD.scala 39:27]
  assign _T_40 = _T_37 | _T_39; // @[LZD.scala 39:25]
  assign _T_41 = {_T_36,_T_40}; // @[Cat.scala 29:58]
  assign _T_42 = _T_34[1:0]; // @[LZD.scala 44:32]
  assign _T_43 = _T_42 != 2'h0; // @[LZD.scala 39:14]
  assign _T_44 = _T_42[1]; // @[LZD.scala 39:21]
  assign _T_45 = _T_42[0]; // @[LZD.scala 39:30]
  assign _T_46 = ~ _T_45; // @[LZD.scala 39:27]
  assign _T_47 = _T_44 | _T_46; // @[LZD.scala 39:25]
  assign _T_48 = {_T_43,_T_47}; // @[Cat.scala 29:58]
  assign _T_49 = _T_41[1]; // @[Shift.scala 12:21]
  assign _T_50 = _T_48[1]; // @[Shift.scala 12:21]
  assign _T_51 = _T_49 | _T_50; // @[LZD.scala 49:16]
  assign _T_52 = ~ _T_50; // @[LZD.scala 49:27]
  assign _T_53 = _T_49 | _T_52; // @[LZD.scala 49:25]
  assign _T_54 = _T_41[0:0]; // @[LZD.scala 49:47]
  assign _T_55 = _T_48[0:0]; // @[LZD.scala 49:59]
  assign _T_56 = _T_49 ? _T_54 : _T_55; // @[LZD.scala 49:35]
  assign _T_58 = {_T_51,_T_53,_T_56}; // @[Cat.scala 29:58]
  assign _T_59 = _T_33[2]; // @[Shift.scala 12:21]
  assign _T_60 = _T_58[2]; // @[Shift.scala 12:21]
  assign _T_61 = _T_59 | _T_60; // @[LZD.scala 49:16]
  assign _T_62 = ~ _T_60; // @[LZD.scala 49:27]
  assign _T_63 = _T_59 | _T_62; // @[LZD.scala 49:25]
  assign _T_64 = _T_33[1:0]; // @[LZD.scala 49:47]
  assign _T_65 = _T_58[1:0]; // @[LZD.scala 49:59]
  assign _T_66 = _T_59 ? _T_64 : _T_65; // @[LZD.scala 49:35]
  assign _T_68 = {_T_61,_T_63,_T_66}; // @[Cat.scala 29:58]
  assign _T_69 = _T_7[7:0]; // @[LZD.scala 44:32]
  assign _T_70 = _T_69[7:4]; // @[LZD.scala 43:32]
  assign _T_71 = _T_70[3:2]; // @[LZD.scala 43:32]
  assign _T_72 = _T_71 != 2'h0; // @[LZD.scala 39:14]
  assign _T_73 = _T_71[1]; // @[LZD.scala 39:21]
  assign _T_74 = _T_71[0]; // @[LZD.scala 39:30]
  assign _T_75 = ~ _T_74; // @[LZD.scala 39:27]
  assign _T_76 = _T_73 | _T_75; // @[LZD.scala 39:25]
  assign _T_77 = {_T_72,_T_76}; // @[Cat.scala 29:58]
  assign _T_78 = _T_70[1:0]; // @[LZD.scala 44:32]
  assign _T_79 = _T_78 != 2'h0; // @[LZD.scala 39:14]
  assign _T_80 = _T_78[1]; // @[LZD.scala 39:21]
  assign _T_81 = _T_78[0]; // @[LZD.scala 39:30]
  assign _T_82 = ~ _T_81; // @[LZD.scala 39:27]
  assign _T_83 = _T_80 | _T_82; // @[LZD.scala 39:25]
  assign _T_84 = {_T_79,_T_83}; // @[Cat.scala 29:58]
  assign _T_85 = _T_77[1]; // @[Shift.scala 12:21]
  assign _T_86 = _T_84[1]; // @[Shift.scala 12:21]
  assign _T_87 = _T_85 | _T_86; // @[LZD.scala 49:16]
  assign _T_88 = ~ _T_86; // @[LZD.scala 49:27]
  assign _T_89 = _T_85 | _T_88; // @[LZD.scala 49:25]
  assign _T_90 = _T_77[0:0]; // @[LZD.scala 49:47]
  assign _T_91 = _T_84[0:0]; // @[LZD.scala 49:59]
  assign _T_92 = _T_85 ? _T_90 : _T_91; // @[LZD.scala 49:35]
  assign _T_94 = {_T_87,_T_89,_T_92}; // @[Cat.scala 29:58]
  assign _T_95 = _T_69[3:0]; // @[LZD.scala 44:32]
  assign _T_96 = _T_95[3:2]; // @[LZD.scala 43:32]
  assign _T_97 = _T_96 != 2'h0; // @[LZD.scala 39:14]
  assign _T_98 = _T_96[1]; // @[LZD.scala 39:21]
  assign _T_99 = _T_96[0]; // @[LZD.scala 39:30]
  assign _T_100 = ~ _T_99; // @[LZD.scala 39:27]
  assign _T_101 = _T_98 | _T_100; // @[LZD.scala 39:25]
  assign _T_102 = {_T_97,_T_101}; // @[Cat.scala 29:58]
  assign _T_103 = _T_95[1:0]; // @[LZD.scala 44:32]
  assign _T_104 = _T_103 != 2'h0; // @[LZD.scala 39:14]
  assign _T_105 = _T_103[1]; // @[LZD.scala 39:21]
  assign _T_106 = _T_103[0]; // @[LZD.scala 39:30]
  assign _T_107 = ~ _T_106; // @[LZD.scala 39:27]
  assign _T_108 = _T_105 | _T_107; // @[LZD.scala 39:25]
  assign _T_109 = {_T_104,_T_108}; // @[Cat.scala 29:58]
  assign _T_110 = _T_102[1]; // @[Shift.scala 12:21]
  assign _T_111 = _T_109[1]; // @[Shift.scala 12:21]
  assign _T_112 = _T_110 | _T_111; // @[LZD.scala 49:16]
  assign _T_113 = ~ _T_111; // @[LZD.scala 49:27]
  assign _T_114 = _T_110 | _T_113; // @[LZD.scala 49:25]
  assign _T_115 = _T_102[0:0]; // @[LZD.scala 49:47]
  assign _T_116 = _T_109[0:0]; // @[LZD.scala 49:59]
  assign _T_117 = _T_110 ? _T_115 : _T_116; // @[LZD.scala 49:35]
  assign _T_119 = {_T_112,_T_114,_T_117}; // @[Cat.scala 29:58]
  assign _T_120 = _T_94[2]; // @[Shift.scala 12:21]
  assign _T_121 = _T_119[2]; // @[Shift.scala 12:21]
  assign _T_122 = _T_120 | _T_121; // @[LZD.scala 49:16]
  assign _T_123 = ~ _T_121; // @[LZD.scala 49:27]
  assign _T_124 = _T_120 | _T_123; // @[LZD.scala 49:25]
  assign _T_125 = _T_94[1:0]; // @[LZD.scala 49:47]
  assign _T_126 = _T_119[1:0]; // @[LZD.scala 49:59]
  assign _T_127 = _T_120 ? _T_125 : _T_126; // @[LZD.scala 49:35]
  assign _T_129 = {_T_122,_T_124,_T_127}; // @[Cat.scala 29:58]
  assign _T_130 = _T_68[3]; // @[Shift.scala 12:21]
  assign _T_131 = _T_129[3]; // @[Shift.scala 12:21]
  assign _T_132 = _T_130 | _T_131; // @[LZD.scala 49:16]
  assign _T_133 = ~ _T_131; // @[LZD.scala 49:27]
  assign _T_134 = _T_130 | _T_133; // @[LZD.scala 49:25]
  assign _T_135 = _T_68[2:0]; // @[LZD.scala 49:47]
  assign _T_136 = _T_129[2:0]; // @[LZD.scala 49:59]
  assign _T_137 = _T_130 ? _T_135 : _T_136; // @[LZD.scala 49:35]
  assign _T_139 = {_T_132,_T_134,_T_137}; // @[Cat.scala 29:58]
  assign _T_140 = _T_6[9:0]; // @[LZD.scala 44:32]
  assign _T_141 = _T_140[9:2]; // @[LZD.scala 43:32]
  assign _T_142 = _T_141[7:4]; // @[LZD.scala 43:32]
  assign _T_143 = _T_142[3:2]; // @[LZD.scala 43:32]
  assign _T_144 = _T_143 != 2'h0; // @[LZD.scala 39:14]
  assign _T_145 = _T_143[1]; // @[LZD.scala 39:21]
  assign _T_146 = _T_143[0]; // @[LZD.scala 39:30]
  assign _T_147 = ~ _T_146; // @[LZD.scala 39:27]
  assign _T_148 = _T_145 | _T_147; // @[LZD.scala 39:25]
  assign _T_149 = {_T_144,_T_148}; // @[Cat.scala 29:58]
  assign _T_150 = _T_142[1:0]; // @[LZD.scala 44:32]
  assign _T_151 = _T_150 != 2'h0; // @[LZD.scala 39:14]
  assign _T_152 = _T_150[1]; // @[LZD.scala 39:21]
  assign _T_153 = _T_150[0]; // @[LZD.scala 39:30]
  assign _T_154 = ~ _T_153; // @[LZD.scala 39:27]
  assign _T_155 = _T_152 | _T_154; // @[LZD.scala 39:25]
  assign _T_156 = {_T_151,_T_155}; // @[Cat.scala 29:58]
  assign _T_157 = _T_149[1]; // @[Shift.scala 12:21]
  assign _T_158 = _T_156[1]; // @[Shift.scala 12:21]
  assign _T_159 = _T_157 | _T_158; // @[LZD.scala 49:16]
  assign _T_160 = ~ _T_158; // @[LZD.scala 49:27]
  assign _T_161 = _T_157 | _T_160; // @[LZD.scala 49:25]
  assign _T_162 = _T_149[0:0]; // @[LZD.scala 49:47]
  assign _T_163 = _T_156[0:0]; // @[LZD.scala 49:59]
  assign _T_164 = _T_157 ? _T_162 : _T_163; // @[LZD.scala 49:35]
  assign _T_166 = {_T_159,_T_161,_T_164}; // @[Cat.scala 29:58]
  assign _T_167 = _T_141[3:0]; // @[LZD.scala 44:32]
  assign _T_168 = _T_167[3:2]; // @[LZD.scala 43:32]
  assign _T_169 = _T_168 != 2'h0; // @[LZD.scala 39:14]
  assign _T_170 = _T_168[1]; // @[LZD.scala 39:21]
  assign _T_171 = _T_168[0]; // @[LZD.scala 39:30]
  assign _T_172 = ~ _T_171; // @[LZD.scala 39:27]
  assign _T_173 = _T_170 | _T_172; // @[LZD.scala 39:25]
  assign _T_174 = {_T_169,_T_173}; // @[Cat.scala 29:58]
  assign _T_175 = _T_167[1:0]; // @[LZD.scala 44:32]
  assign _T_176 = _T_175 != 2'h0; // @[LZD.scala 39:14]
  assign _T_177 = _T_175[1]; // @[LZD.scala 39:21]
  assign _T_178 = _T_175[0]; // @[LZD.scala 39:30]
  assign _T_179 = ~ _T_178; // @[LZD.scala 39:27]
  assign _T_180 = _T_177 | _T_179; // @[LZD.scala 39:25]
  assign _T_181 = {_T_176,_T_180}; // @[Cat.scala 29:58]
  assign _T_182 = _T_174[1]; // @[Shift.scala 12:21]
  assign _T_183 = _T_181[1]; // @[Shift.scala 12:21]
  assign _T_184 = _T_182 | _T_183; // @[LZD.scala 49:16]
  assign _T_185 = ~ _T_183; // @[LZD.scala 49:27]
  assign _T_186 = _T_182 | _T_185; // @[LZD.scala 49:25]
  assign _T_187 = _T_174[0:0]; // @[LZD.scala 49:47]
  assign _T_188 = _T_181[0:0]; // @[LZD.scala 49:59]
  assign _T_189 = _T_182 ? _T_187 : _T_188; // @[LZD.scala 49:35]
  assign _T_191 = {_T_184,_T_186,_T_189}; // @[Cat.scala 29:58]
  assign _T_192 = _T_166[2]; // @[Shift.scala 12:21]
  assign _T_193 = _T_191[2]; // @[Shift.scala 12:21]
  assign _T_194 = _T_192 | _T_193; // @[LZD.scala 49:16]
  assign _T_195 = ~ _T_193; // @[LZD.scala 49:27]
  assign _T_196 = _T_192 | _T_195; // @[LZD.scala 49:25]
  assign _T_197 = _T_166[1:0]; // @[LZD.scala 49:47]
  assign _T_198 = _T_191[1:0]; // @[LZD.scala 49:59]
  assign _T_199 = _T_192 ? _T_197 : _T_198; // @[LZD.scala 49:35]
  assign _T_201 = {_T_194,_T_196,_T_199}; // @[Cat.scala 29:58]
  assign _T_202 = _T_140[1:0]; // @[LZD.scala 44:32]
  assign _T_203 = _T_202 != 2'h0; // @[LZD.scala 39:14]
  assign _T_204 = _T_202[1]; // @[LZD.scala 39:21]
  assign _T_205 = _T_202[0]; // @[LZD.scala 39:30]
  assign _T_206 = ~ _T_205; // @[LZD.scala 39:27]
  assign _T_207 = _T_204 | _T_206; // @[LZD.scala 39:25]
  assign _T_209 = _T_201[3]; // @[Shift.scala 12:21]
  assign _T_211 = {1'h1,_T_203,_T_207}; // @[Cat.scala 29:58]
  assign _T_212 = _T_201[2:0]; // @[LZD.scala 55:32]
  assign _T_213 = _T_209 ? _T_212 : _T_211; // @[LZD.scala 55:20]
  assign _T_214 = {_T_209,_T_213}; // @[Cat.scala 29:58]
  assign _T_215 = _T_139[4]; // @[Shift.scala 12:21]
  assign _T_217 = _T_139[3:0]; // @[LZD.scala 55:32]
  assign _T_218 = _T_215 ? _T_217 : _T_214; // @[LZD.scala 55:20]
  assign _T_219 = {_T_215,_T_218}; // @[Cat.scala 29:58]
  assign _T_220 = ~ _T_219; // @[convert.scala 21:22]
  assign _T_221 = io_A[24:0]; // @[convert.scala 22:36]
  assign _T_222 = _T_220 < 5'h19; // @[Shift.scala 16:24]
  assign _T_224 = _T_220[4]; // @[Shift.scala 12:21]
  assign _T_225 = _T_221[8:0]; // @[Shift.scala 64:52]
  assign _T_227 = {_T_225,16'h0}; // @[Cat.scala 29:58]
  assign _T_228 = _T_224 ? _T_227 : _T_221; // @[Shift.scala 64:27]
  assign _T_229 = _T_220[3:0]; // @[Shift.scala 66:70]
  assign _T_230 = _T_229[3]; // @[Shift.scala 12:21]
  assign _T_231 = _T_228[16:0]; // @[Shift.scala 64:52]
  assign _T_233 = {_T_231,8'h0}; // @[Cat.scala 29:58]
  assign _T_234 = _T_230 ? _T_233 : _T_228; // @[Shift.scala 64:27]
  assign _T_235 = _T_229[2:0]; // @[Shift.scala 66:70]
  assign _T_236 = _T_235[2]; // @[Shift.scala 12:21]
  assign _T_237 = _T_234[20:0]; // @[Shift.scala 64:52]
  assign _T_239 = {_T_237,4'h0}; // @[Cat.scala 29:58]
  assign _T_240 = _T_236 ? _T_239 : _T_234; // @[Shift.scala 64:27]
  assign _T_241 = _T_235[1:0]; // @[Shift.scala 66:70]
  assign _T_242 = _T_241[1]; // @[Shift.scala 12:21]
  assign _T_243 = _T_240[22:0]; // @[Shift.scala 64:52]
  assign _T_245 = {_T_243,2'h0}; // @[Cat.scala 29:58]
  assign _T_246 = _T_242 ? _T_245 : _T_240; // @[Shift.scala 64:27]
  assign _T_247 = _T_241[0:0]; // @[Shift.scala 66:70]
  assign _T_249 = _T_246[23:0]; // @[Shift.scala 64:52]
  assign _T_250 = {_T_249,1'h0}; // @[Cat.scala 29:58]
  assign _T_251 = _T_247 ? _T_250 : _T_246; // @[Shift.scala 64:27]
  assign _T_252 = _T_222 ? _T_251 : 25'h0; // @[Shift.scala 16:10]
  assign _T_253 = _T_252[24:22]; // @[convert.scala 23:34]
  assign decA_fraction = _T_252[21:0]; // @[convert.scala 24:34]
  assign _T_255 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_257 = _T_3 ? _T_220 : _T_219; // @[convert.scala 25:42]
  assign _T_260 = ~ _T_253; // @[convert.scala 26:67]
  assign _T_261 = _T_1 ? _T_260 : _T_253; // @[convert.scala 26:51]
  assign _T_262 = {_T_255,_T_257,_T_261}; // @[Cat.scala 29:58]
  assign _T_264 = io_A[26:0]; // @[convert.scala 29:56]
  assign _T_265 = _T_264 != 27'h0; // @[convert.scala 29:60]
  assign _T_266 = ~ _T_265; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_266; // @[convert.scala 29:39]
  assign _T_269 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_269 & _T_266; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_262); // @[convert.scala 32:24]
  assign _T_278 = io_B[27]; // @[convert.scala 18:24]
  assign _T_279 = io_B[26]; // @[convert.scala 18:40]
  assign _T_280 = _T_278 ^ _T_279; // @[convert.scala 18:36]
  assign _T_281 = io_B[26:1]; // @[convert.scala 19:24]
  assign _T_282 = io_B[25:0]; // @[convert.scala 19:43]
  assign _T_283 = _T_281 ^ _T_282; // @[convert.scala 19:39]
  assign _T_284 = _T_283[25:10]; // @[LZD.scala 43:32]
  assign _T_285 = _T_284[15:8]; // @[LZD.scala 43:32]
  assign _T_286 = _T_285[7:4]; // @[LZD.scala 43:32]
  assign _T_287 = _T_286[3:2]; // @[LZD.scala 43:32]
  assign _T_288 = _T_287 != 2'h0; // @[LZD.scala 39:14]
  assign _T_289 = _T_287[1]; // @[LZD.scala 39:21]
  assign _T_290 = _T_287[0]; // @[LZD.scala 39:30]
  assign _T_291 = ~ _T_290; // @[LZD.scala 39:27]
  assign _T_292 = _T_289 | _T_291; // @[LZD.scala 39:25]
  assign _T_293 = {_T_288,_T_292}; // @[Cat.scala 29:58]
  assign _T_294 = _T_286[1:0]; // @[LZD.scala 44:32]
  assign _T_295 = _T_294 != 2'h0; // @[LZD.scala 39:14]
  assign _T_296 = _T_294[1]; // @[LZD.scala 39:21]
  assign _T_297 = _T_294[0]; // @[LZD.scala 39:30]
  assign _T_298 = ~ _T_297; // @[LZD.scala 39:27]
  assign _T_299 = _T_296 | _T_298; // @[LZD.scala 39:25]
  assign _T_300 = {_T_295,_T_299}; // @[Cat.scala 29:58]
  assign _T_301 = _T_293[1]; // @[Shift.scala 12:21]
  assign _T_302 = _T_300[1]; // @[Shift.scala 12:21]
  assign _T_303 = _T_301 | _T_302; // @[LZD.scala 49:16]
  assign _T_304 = ~ _T_302; // @[LZD.scala 49:27]
  assign _T_305 = _T_301 | _T_304; // @[LZD.scala 49:25]
  assign _T_306 = _T_293[0:0]; // @[LZD.scala 49:47]
  assign _T_307 = _T_300[0:0]; // @[LZD.scala 49:59]
  assign _T_308 = _T_301 ? _T_306 : _T_307; // @[LZD.scala 49:35]
  assign _T_310 = {_T_303,_T_305,_T_308}; // @[Cat.scala 29:58]
  assign _T_311 = _T_285[3:0]; // @[LZD.scala 44:32]
  assign _T_312 = _T_311[3:2]; // @[LZD.scala 43:32]
  assign _T_313 = _T_312 != 2'h0; // @[LZD.scala 39:14]
  assign _T_314 = _T_312[1]; // @[LZD.scala 39:21]
  assign _T_315 = _T_312[0]; // @[LZD.scala 39:30]
  assign _T_316 = ~ _T_315; // @[LZD.scala 39:27]
  assign _T_317 = _T_314 | _T_316; // @[LZD.scala 39:25]
  assign _T_318 = {_T_313,_T_317}; // @[Cat.scala 29:58]
  assign _T_319 = _T_311[1:0]; // @[LZD.scala 44:32]
  assign _T_320 = _T_319 != 2'h0; // @[LZD.scala 39:14]
  assign _T_321 = _T_319[1]; // @[LZD.scala 39:21]
  assign _T_322 = _T_319[0]; // @[LZD.scala 39:30]
  assign _T_323 = ~ _T_322; // @[LZD.scala 39:27]
  assign _T_324 = _T_321 | _T_323; // @[LZD.scala 39:25]
  assign _T_325 = {_T_320,_T_324}; // @[Cat.scala 29:58]
  assign _T_326 = _T_318[1]; // @[Shift.scala 12:21]
  assign _T_327 = _T_325[1]; // @[Shift.scala 12:21]
  assign _T_328 = _T_326 | _T_327; // @[LZD.scala 49:16]
  assign _T_329 = ~ _T_327; // @[LZD.scala 49:27]
  assign _T_330 = _T_326 | _T_329; // @[LZD.scala 49:25]
  assign _T_331 = _T_318[0:0]; // @[LZD.scala 49:47]
  assign _T_332 = _T_325[0:0]; // @[LZD.scala 49:59]
  assign _T_333 = _T_326 ? _T_331 : _T_332; // @[LZD.scala 49:35]
  assign _T_335 = {_T_328,_T_330,_T_333}; // @[Cat.scala 29:58]
  assign _T_336 = _T_310[2]; // @[Shift.scala 12:21]
  assign _T_337 = _T_335[2]; // @[Shift.scala 12:21]
  assign _T_338 = _T_336 | _T_337; // @[LZD.scala 49:16]
  assign _T_339 = ~ _T_337; // @[LZD.scala 49:27]
  assign _T_340 = _T_336 | _T_339; // @[LZD.scala 49:25]
  assign _T_341 = _T_310[1:0]; // @[LZD.scala 49:47]
  assign _T_342 = _T_335[1:0]; // @[LZD.scala 49:59]
  assign _T_343 = _T_336 ? _T_341 : _T_342; // @[LZD.scala 49:35]
  assign _T_345 = {_T_338,_T_340,_T_343}; // @[Cat.scala 29:58]
  assign _T_346 = _T_284[7:0]; // @[LZD.scala 44:32]
  assign _T_347 = _T_346[7:4]; // @[LZD.scala 43:32]
  assign _T_348 = _T_347[3:2]; // @[LZD.scala 43:32]
  assign _T_349 = _T_348 != 2'h0; // @[LZD.scala 39:14]
  assign _T_350 = _T_348[1]; // @[LZD.scala 39:21]
  assign _T_351 = _T_348[0]; // @[LZD.scala 39:30]
  assign _T_352 = ~ _T_351; // @[LZD.scala 39:27]
  assign _T_353 = _T_350 | _T_352; // @[LZD.scala 39:25]
  assign _T_354 = {_T_349,_T_353}; // @[Cat.scala 29:58]
  assign _T_355 = _T_347[1:0]; // @[LZD.scala 44:32]
  assign _T_356 = _T_355 != 2'h0; // @[LZD.scala 39:14]
  assign _T_357 = _T_355[1]; // @[LZD.scala 39:21]
  assign _T_358 = _T_355[0]; // @[LZD.scala 39:30]
  assign _T_359 = ~ _T_358; // @[LZD.scala 39:27]
  assign _T_360 = _T_357 | _T_359; // @[LZD.scala 39:25]
  assign _T_361 = {_T_356,_T_360}; // @[Cat.scala 29:58]
  assign _T_362 = _T_354[1]; // @[Shift.scala 12:21]
  assign _T_363 = _T_361[1]; // @[Shift.scala 12:21]
  assign _T_364 = _T_362 | _T_363; // @[LZD.scala 49:16]
  assign _T_365 = ~ _T_363; // @[LZD.scala 49:27]
  assign _T_366 = _T_362 | _T_365; // @[LZD.scala 49:25]
  assign _T_367 = _T_354[0:0]; // @[LZD.scala 49:47]
  assign _T_368 = _T_361[0:0]; // @[LZD.scala 49:59]
  assign _T_369 = _T_362 ? _T_367 : _T_368; // @[LZD.scala 49:35]
  assign _T_371 = {_T_364,_T_366,_T_369}; // @[Cat.scala 29:58]
  assign _T_372 = _T_346[3:0]; // @[LZD.scala 44:32]
  assign _T_373 = _T_372[3:2]; // @[LZD.scala 43:32]
  assign _T_374 = _T_373 != 2'h0; // @[LZD.scala 39:14]
  assign _T_375 = _T_373[1]; // @[LZD.scala 39:21]
  assign _T_376 = _T_373[0]; // @[LZD.scala 39:30]
  assign _T_377 = ~ _T_376; // @[LZD.scala 39:27]
  assign _T_378 = _T_375 | _T_377; // @[LZD.scala 39:25]
  assign _T_379 = {_T_374,_T_378}; // @[Cat.scala 29:58]
  assign _T_380 = _T_372[1:0]; // @[LZD.scala 44:32]
  assign _T_381 = _T_380 != 2'h0; // @[LZD.scala 39:14]
  assign _T_382 = _T_380[1]; // @[LZD.scala 39:21]
  assign _T_383 = _T_380[0]; // @[LZD.scala 39:30]
  assign _T_384 = ~ _T_383; // @[LZD.scala 39:27]
  assign _T_385 = _T_382 | _T_384; // @[LZD.scala 39:25]
  assign _T_386 = {_T_381,_T_385}; // @[Cat.scala 29:58]
  assign _T_387 = _T_379[1]; // @[Shift.scala 12:21]
  assign _T_388 = _T_386[1]; // @[Shift.scala 12:21]
  assign _T_389 = _T_387 | _T_388; // @[LZD.scala 49:16]
  assign _T_390 = ~ _T_388; // @[LZD.scala 49:27]
  assign _T_391 = _T_387 | _T_390; // @[LZD.scala 49:25]
  assign _T_392 = _T_379[0:0]; // @[LZD.scala 49:47]
  assign _T_393 = _T_386[0:0]; // @[LZD.scala 49:59]
  assign _T_394 = _T_387 ? _T_392 : _T_393; // @[LZD.scala 49:35]
  assign _T_396 = {_T_389,_T_391,_T_394}; // @[Cat.scala 29:58]
  assign _T_397 = _T_371[2]; // @[Shift.scala 12:21]
  assign _T_398 = _T_396[2]; // @[Shift.scala 12:21]
  assign _T_399 = _T_397 | _T_398; // @[LZD.scala 49:16]
  assign _T_400 = ~ _T_398; // @[LZD.scala 49:27]
  assign _T_401 = _T_397 | _T_400; // @[LZD.scala 49:25]
  assign _T_402 = _T_371[1:0]; // @[LZD.scala 49:47]
  assign _T_403 = _T_396[1:0]; // @[LZD.scala 49:59]
  assign _T_404 = _T_397 ? _T_402 : _T_403; // @[LZD.scala 49:35]
  assign _T_406 = {_T_399,_T_401,_T_404}; // @[Cat.scala 29:58]
  assign _T_407 = _T_345[3]; // @[Shift.scala 12:21]
  assign _T_408 = _T_406[3]; // @[Shift.scala 12:21]
  assign _T_409 = _T_407 | _T_408; // @[LZD.scala 49:16]
  assign _T_410 = ~ _T_408; // @[LZD.scala 49:27]
  assign _T_411 = _T_407 | _T_410; // @[LZD.scala 49:25]
  assign _T_412 = _T_345[2:0]; // @[LZD.scala 49:47]
  assign _T_413 = _T_406[2:0]; // @[LZD.scala 49:59]
  assign _T_414 = _T_407 ? _T_412 : _T_413; // @[LZD.scala 49:35]
  assign _T_416 = {_T_409,_T_411,_T_414}; // @[Cat.scala 29:58]
  assign _T_417 = _T_283[9:0]; // @[LZD.scala 44:32]
  assign _T_418 = _T_417[9:2]; // @[LZD.scala 43:32]
  assign _T_419 = _T_418[7:4]; // @[LZD.scala 43:32]
  assign _T_420 = _T_419[3:2]; // @[LZD.scala 43:32]
  assign _T_421 = _T_420 != 2'h0; // @[LZD.scala 39:14]
  assign _T_422 = _T_420[1]; // @[LZD.scala 39:21]
  assign _T_423 = _T_420[0]; // @[LZD.scala 39:30]
  assign _T_424 = ~ _T_423; // @[LZD.scala 39:27]
  assign _T_425 = _T_422 | _T_424; // @[LZD.scala 39:25]
  assign _T_426 = {_T_421,_T_425}; // @[Cat.scala 29:58]
  assign _T_427 = _T_419[1:0]; // @[LZD.scala 44:32]
  assign _T_428 = _T_427 != 2'h0; // @[LZD.scala 39:14]
  assign _T_429 = _T_427[1]; // @[LZD.scala 39:21]
  assign _T_430 = _T_427[0]; // @[LZD.scala 39:30]
  assign _T_431 = ~ _T_430; // @[LZD.scala 39:27]
  assign _T_432 = _T_429 | _T_431; // @[LZD.scala 39:25]
  assign _T_433 = {_T_428,_T_432}; // @[Cat.scala 29:58]
  assign _T_434 = _T_426[1]; // @[Shift.scala 12:21]
  assign _T_435 = _T_433[1]; // @[Shift.scala 12:21]
  assign _T_436 = _T_434 | _T_435; // @[LZD.scala 49:16]
  assign _T_437 = ~ _T_435; // @[LZD.scala 49:27]
  assign _T_438 = _T_434 | _T_437; // @[LZD.scala 49:25]
  assign _T_439 = _T_426[0:0]; // @[LZD.scala 49:47]
  assign _T_440 = _T_433[0:0]; // @[LZD.scala 49:59]
  assign _T_441 = _T_434 ? _T_439 : _T_440; // @[LZD.scala 49:35]
  assign _T_443 = {_T_436,_T_438,_T_441}; // @[Cat.scala 29:58]
  assign _T_444 = _T_418[3:0]; // @[LZD.scala 44:32]
  assign _T_445 = _T_444[3:2]; // @[LZD.scala 43:32]
  assign _T_446 = _T_445 != 2'h0; // @[LZD.scala 39:14]
  assign _T_447 = _T_445[1]; // @[LZD.scala 39:21]
  assign _T_448 = _T_445[0]; // @[LZD.scala 39:30]
  assign _T_449 = ~ _T_448; // @[LZD.scala 39:27]
  assign _T_450 = _T_447 | _T_449; // @[LZD.scala 39:25]
  assign _T_451 = {_T_446,_T_450}; // @[Cat.scala 29:58]
  assign _T_452 = _T_444[1:0]; // @[LZD.scala 44:32]
  assign _T_453 = _T_452 != 2'h0; // @[LZD.scala 39:14]
  assign _T_454 = _T_452[1]; // @[LZD.scala 39:21]
  assign _T_455 = _T_452[0]; // @[LZD.scala 39:30]
  assign _T_456 = ~ _T_455; // @[LZD.scala 39:27]
  assign _T_457 = _T_454 | _T_456; // @[LZD.scala 39:25]
  assign _T_458 = {_T_453,_T_457}; // @[Cat.scala 29:58]
  assign _T_459 = _T_451[1]; // @[Shift.scala 12:21]
  assign _T_460 = _T_458[1]; // @[Shift.scala 12:21]
  assign _T_461 = _T_459 | _T_460; // @[LZD.scala 49:16]
  assign _T_462 = ~ _T_460; // @[LZD.scala 49:27]
  assign _T_463 = _T_459 | _T_462; // @[LZD.scala 49:25]
  assign _T_464 = _T_451[0:0]; // @[LZD.scala 49:47]
  assign _T_465 = _T_458[0:0]; // @[LZD.scala 49:59]
  assign _T_466 = _T_459 ? _T_464 : _T_465; // @[LZD.scala 49:35]
  assign _T_468 = {_T_461,_T_463,_T_466}; // @[Cat.scala 29:58]
  assign _T_469 = _T_443[2]; // @[Shift.scala 12:21]
  assign _T_470 = _T_468[2]; // @[Shift.scala 12:21]
  assign _T_471 = _T_469 | _T_470; // @[LZD.scala 49:16]
  assign _T_472 = ~ _T_470; // @[LZD.scala 49:27]
  assign _T_473 = _T_469 | _T_472; // @[LZD.scala 49:25]
  assign _T_474 = _T_443[1:0]; // @[LZD.scala 49:47]
  assign _T_475 = _T_468[1:0]; // @[LZD.scala 49:59]
  assign _T_476 = _T_469 ? _T_474 : _T_475; // @[LZD.scala 49:35]
  assign _T_478 = {_T_471,_T_473,_T_476}; // @[Cat.scala 29:58]
  assign _T_479 = _T_417[1:0]; // @[LZD.scala 44:32]
  assign _T_480 = _T_479 != 2'h0; // @[LZD.scala 39:14]
  assign _T_481 = _T_479[1]; // @[LZD.scala 39:21]
  assign _T_482 = _T_479[0]; // @[LZD.scala 39:30]
  assign _T_483 = ~ _T_482; // @[LZD.scala 39:27]
  assign _T_484 = _T_481 | _T_483; // @[LZD.scala 39:25]
  assign _T_486 = _T_478[3]; // @[Shift.scala 12:21]
  assign _T_488 = {1'h1,_T_480,_T_484}; // @[Cat.scala 29:58]
  assign _T_489 = _T_478[2:0]; // @[LZD.scala 55:32]
  assign _T_490 = _T_486 ? _T_489 : _T_488; // @[LZD.scala 55:20]
  assign _T_491 = {_T_486,_T_490}; // @[Cat.scala 29:58]
  assign _T_492 = _T_416[4]; // @[Shift.scala 12:21]
  assign _T_494 = _T_416[3:0]; // @[LZD.scala 55:32]
  assign _T_495 = _T_492 ? _T_494 : _T_491; // @[LZD.scala 55:20]
  assign _T_496 = {_T_492,_T_495}; // @[Cat.scala 29:58]
  assign _T_497 = ~ _T_496; // @[convert.scala 21:22]
  assign _T_498 = io_B[24:0]; // @[convert.scala 22:36]
  assign _T_499 = _T_497 < 5'h19; // @[Shift.scala 16:24]
  assign _T_501 = _T_497[4]; // @[Shift.scala 12:21]
  assign _T_502 = _T_498[8:0]; // @[Shift.scala 64:52]
  assign _T_504 = {_T_502,16'h0}; // @[Cat.scala 29:58]
  assign _T_505 = _T_501 ? _T_504 : _T_498; // @[Shift.scala 64:27]
  assign _T_506 = _T_497[3:0]; // @[Shift.scala 66:70]
  assign _T_507 = _T_506[3]; // @[Shift.scala 12:21]
  assign _T_508 = _T_505[16:0]; // @[Shift.scala 64:52]
  assign _T_510 = {_T_508,8'h0}; // @[Cat.scala 29:58]
  assign _T_511 = _T_507 ? _T_510 : _T_505; // @[Shift.scala 64:27]
  assign _T_512 = _T_506[2:0]; // @[Shift.scala 66:70]
  assign _T_513 = _T_512[2]; // @[Shift.scala 12:21]
  assign _T_514 = _T_511[20:0]; // @[Shift.scala 64:52]
  assign _T_516 = {_T_514,4'h0}; // @[Cat.scala 29:58]
  assign _T_517 = _T_513 ? _T_516 : _T_511; // @[Shift.scala 64:27]
  assign _T_518 = _T_512[1:0]; // @[Shift.scala 66:70]
  assign _T_519 = _T_518[1]; // @[Shift.scala 12:21]
  assign _T_520 = _T_517[22:0]; // @[Shift.scala 64:52]
  assign _T_522 = {_T_520,2'h0}; // @[Cat.scala 29:58]
  assign _T_523 = _T_519 ? _T_522 : _T_517; // @[Shift.scala 64:27]
  assign _T_524 = _T_518[0:0]; // @[Shift.scala 66:70]
  assign _T_526 = _T_523[23:0]; // @[Shift.scala 64:52]
  assign _T_527 = {_T_526,1'h0}; // @[Cat.scala 29:58]
  assign _T_528 = _T_524 ? _T_527 : _T_523; // @[Shift.scala 64:27]
  assign _T_529 = _T_499 ? _T_528 : 25'h0; // @[Shift.scala 16:10]
  assign _T_530 = _T_529[24:22]; // @[convert.scala 23:34]
  assign decB_fraction = _T_529[21:0]; // @[convert.scala 24:34]
  assign _T_532 = _T_280 == 1'h0; // @[convert.scala 25:26]
  assign _T_534 = _T_280 ? _T_497 : _T_496; // @[convert.scala 25:42]
  assign _T_537 = ~ _T_530; // @[convert.scala 26:67]
  assign _T_538 = _T_278 ? _T_537 : _T_530; // @[convert.scala 26:51]
  assign _T_539 = {_T_532,_T_534,_T_538}; // @[Cat.scala 29:58]
  assign _T_541 = io_B[26:0]; // @[convert.scala 29:56]
  assign _T_542 = _T_541 != 27'h0; // @[convert.scala 29:60]
  assign _T_543 = ~ _T_542; // @[convert.scala 29:41]
  assign decB_isNaR = _T_278 & _T_543; // @[convert.scala 29:39]
  assign _T_546 = _T_278 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_546 & _T_543; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_539); // @[convert.scala 32:24]
  assign _T_554 = ~ _T_1; // @[PositMultiplier.scala 43:34]
  assign _T_556 = {_T_1,_T_554,decA_fraction}; // @[Cat.scala 29:58]
  assign sigA = $signed(_T_556); // @[PositMultiplier.scala 43:61]
  assign _T_557 = ~ _T_278; // @[PositMultiplier.scala 44:34]
  assign _T_559 = {_T_278,_T_557,decB_fraction}; // @[Cat.scala 29:58]
  assign sigB = $signed(_T_559); // @[PositMultiplier.scala 44:61]
  assign _T_560 = $signed(sigA) * $signed(sigB); // @[PositMultiplier.scala 45:25]
  assign sigP = $unsigned(_T_560); // @[PositMultiplier.scala 45:33]
  assign head2 = sigP[47:46]; // @[PositMultiplier.scala 46:28]
  assign _T_561 = head2[1]; // @[PositMultiplier.scala 47:31]
  assign _T_562 = ~ _T_561; // @[PositMultiplier.scala 47:25]
  assign _T_563 = head2[0]; // @[PositMultiplier.scala 47:42]
  assign addTwo = _T_562 & _T_563; // @[PositMultiplier.scala 47:35]
  assign _T_564 = sigP[47]; // @[PositMultiplier.scala 49:23]
  assign _T_565 = sigP[45]; // @[PositMultiplier.scala 49:49]
  assign addOne = _T_564 ^ _T_565; // @[PositMultiplier.scala 49:43]
  assign _T_566 = {addTwo,addOne}; // @[Cat.scala 29:58]
  assign expBias = {1'b0,$signed(_T_566)}; // @[PositMultiplier.scala 50:39]
  assign _T_567 = sigP[44:0]; // @[PositMultiplier.scala 53:81]
  assign _T_568 = sigP[43:0]; // @[PositMultiplier.scala 54:81]
  assign _T_569 = {_T_568, 1'h0}; // @[PositMultiplier.scala 54:104]
  assign frac = addOne ? _T_567 : _T_569; // @[PositMultiplier.scala 51:22]
  assign _T_570 = $signed(decA_scale) + $signed(decB_scale); // @[PositMultiplier.scala 56:30]
  assign _GEN_0 = {{7{expBias[2]}},expBias}; // @[PositMultiplier.scala 56:44]
  assign _T_572 = $signed(_T_570) + $signed(_GEN_0); // @[PositMultiplier.scala 56:44]
  assign mulScale = $signed(_T_572); // @[PositMultiplier.scala 56:44]
  assign underflow = $signed(mulScale) < $signed(-10'shd1); // @[PositMultiplier.scala 57:28]
  assign overflow = $signed(mulScale) > $signed(10'shd0); // @[PositMultiplier.scala 58:28]
  assign decM_sign = sigP[47:47]; // @[PositMultiplier.scala 62:29]
  assign _T_575 = underflow ? $signed(-10'shd1) : $signed(mulScale); // @[Mux.scala 87:16]
  assign _T_576 = overflow ? $signed(10'shd0) : $signed(_T_575); // @[Mux.scala 87:16]
  assign decM_fraction = frac[44:23]; // @[PositMultiplier.scala 70:29]
  assign decM_isNaR = decA_isNaR | decB_isNaR; // @[PositMultiplier.scala 71:31]
  assign decM_isZero = decA_isZero | decB_isZero; // @[PositMultiplier.scala 72:32]
  assign grsTmp = frac[22:0]; // @[PositMultiplier.scala 75:30]
  assign _T_580 = grsTmp[22:21]; // @[PositMultiplier.scala 78:32]
  assign _T_581 = grsTmp[20:0]; // @[PositMultiplier.scala 78:48]
  assign _T_582 = _T_581 != 21'h0; // @[PositMultiplier.scala 78:52]
  assign _GEN_1 = _T_576[8:0]; // @[PositMultiplier.scala 60:23 PositMultiplier.scala 63:17]
  assign decM_scale = $signed(_GEN_1); // @[PositMultiplier.scala 60:23 PositMultiplier.scala 63:17]
  assign _T_585 = decM_scale[2:0]; // @[convert.scala 46:61]
  assign _T_586 = ~ _T_585; // @[convert.scala 46:52]
  assign _T_588 = decM_sign ? _T_586 : _T_585; // @[convert.scala 46:42]
  assign _T_589 = decM_scale[8:3]; // @[convert.scala 48:34]
  assign _T_590 = _T_589[5:5]; // @[convert.scala 49:36]
  assign _T_592 = ~ _T_589; // @[convert.scala 50:36]
  assign _T_593 = $signed(_T_592); // @[convert.scala 50:36]
  assign _T_594 = _T_590 ? $signed(_T_593) : $signed(_T_589); // @[convert.scala 50:28]
  assign _T_595 = _T_590 ^ decM_sign; // @[convert.scala 51:31]
  assign _T_596 = ~ _T_595; // @[convert.scala 52:43]
  assign _T_600 = {_T_596,_T_595,_T_588,decM_fraction,_T_580,_T_582}; // @[Cat.scala 29:58]
  assign _T_601 = $unsigned(_T_594); // @[Shift.scala 39:17]
  assign _T_602 = _T_601 < 6'h1e; // @[Shift.scala 39:24]
  assign _T_603 = _T_594[4:0]; // @[Shift.scala 40:44]
  assign _T_604 = _T_600[29:16]; // @[Shift.scala 90:30]
  assign _T_605 = _T_600[15:0]; // @[Shift.scala 90:48]
  assign _T_606 = _T_605 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_2 = {{13'd0}, _T_606}; // @[Shift.scala 90:39]
  assign _T_607 = _T_604 | _GEN_2; // @[Shift.scala 90:39]
  assign _T_608 = _T_603[4]; // @[Shift.scala 12:21]
  assign _T_609 = _T_600[29]; // @[Shift.scala 12:21]
  assign _T_611 = _T_609 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_612 = {_T_611,_T_607}; // @[Cat.scala 29:58]
  assign _T_613 = _T_608 ? _T_612 : _T_600; // @[Shift.scala 91:22]
  assign _T_614 = _T_603[3:0]; // @[Shift.scala 92:77]
  assign _T_615 = _T_613[29:8]; // @[Shift.scala 90:30]
  assign _T_616 = _T_613[7:0]; // @[Shift.scala 90:48]
  assign _T_617 = _T_616 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_3 = {{21'd0}, _T_617}; // @[Shift.scala 90:39]
  assign _T_618 = _T_615 | _GEN_3; // @[Shift.scala 90:39]
  assign _T_619 = _T_614[3]; // @[Shift.scala 12:21]
  assign _T_620 = _T_613[29]; // @[Shift.scala 12:21]
  assign _T_622 = _T_620 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_623 = {_T_622,_T_618}; // @[Cat.scala 29:58]
  assign _T_624 = _T_619 ? _T_623 : _T_613; // @[Shift.scala 91:22]
  assign _T_625 = _T_614[2:0]; // @[Shift.scala 92:77]
  assign _T_626 = _T_624[29:4]; // @[Shift.scala 90:30]
  assign _T_627 = _T_624[3:0]; // @[Shift.scala 90:48]
  assign _T_628 = _T_627 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_4 = {{25'd0}, _T_628}; // @[Shift.scala 90:39]
  assign _T_629 = _T_626 | _GEN_4; // @[Shift.scala 90:39]
  assign _T_630 = _T_625[2]; // @[Shift.scala 12:21]
  assign _T_631 = _T_624[29]; // @[Shift.scala 12:21]
  assign _T_633 = _T_631 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_634 = {_T_633,_T_629}; // @[Cat.scala 29:58]
  assign _T_635 = _T_630 ? _T_634 : _T_624; // @[Shift.scala 91:22]
  assign _T_636 = _T_625[1:0]; // @[Shift.scala 92:77]
  assign _T_637 = _T_635[29:2]; // @[Shift.scala 90:30]
  assign _T_638 = _T_635[1:0]; // @[Shift.scala 90:48]
  assign _T_639 = _T_638 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_5 = {{27'd0}, _T_639}; // @[Shift.scala 90:39]
  assign _T_640 = _T_637 | _GEN_5; // @[Shift.scala 90:39]
  assign _T_641 = _T_636[1]; // @[Shift.scala 12:21]
  assign _T_642 = _T_635[29]; // @[Shift.scala 12:21]
  assign _T_644 = _T_642 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_645 = {_T_644,_T_640}; // @[Cat.scala 29:58]
  assign _T_646 = _T_641 ? _T_645 : _T_635; // @[Shift.scala 91:22]
  assign _T_647 = _T_636[0:0]; // @[Shift.scala 92:77]
  assign _T_648 = _T_646[29:1]; // @[Shift.scala 90:30]
  assign _T_649 = _T_646[0:0]; // @[Shift.scala 90:48]
  assign _GEN_6 = {{28'd0}, _T_649}; // @[Shift.scala 90:39]
  assign _T_651 = _T_648 | _GEN_6; // @[Shift.scala 90:39]
  assign _T_653 = _T_646[29]; // @[Shift.scala 12:21]
  assign _T_654 = {_T_653,_T_651}; // @[Cat.scala 29:58]
  assign _T_655 = _T_647 ? _T_654 : _T_646; // @[Shift.scala 91:22]
  assign _T_658 = _T_609 ? 30'h3fffffff : 30'h0; // @[Bitwise.scala 71:12]
  assign _T_659 = _T_602 ? _T_655 : _T_658; // @[Shift.scala 39:10]
  assign _T_660 = _T_659[3]; // @[convert.scala 55:31]
  assign _T_661 = _T_659[2]; // @[convert.scala 56:31]
  assign _T_662 = _T_659[1]; // @[convert.scala 57:31]
  assign _T_663 = _T_659[0]; // @[convert.scala 58:31]
  assign _T_664 = _T_659[29:3]; // @[convert.scala 59:69]
  assign _T_665 = _T_664 != 27'h0; // @[convert.scala 59:81]
  assign _T_666 = ~ _T_665; // @[convert.scala 59:50]
  assign _T_668 = _T_664 == 27'h7ffffff; // @[convert.scala 60:81]
  assign _T_669 = _T_660 | _T_662; // @[convert.scala 61:44]
  assign _T_670 = _T_669 | _T_663; // @[convert.scala 61:52]
  assign _T_671 = _T_661 & _T_670; // @[convert.scala 61:36]
  assign _T_672 = ~ _T_668; // @[convert.scala 62:63]
  assign _T_673 = _T_672 & _T_671; // @[convert.scala 62:103]
  assign _T_674 = _T_666 | _T_673; // @[convert.scala 62:60]
  assign _GEN_7 = {{26'd0}, _T_674}; // @[convert.scala 63:56]
  assign _T_677 = _T_664 + _GEN_7; // @[convert.scala 63:56]
  assign _T_678 = {decM_sign,_T_677}; // @[Cat.scala 29:58]
  assign _T_680 = decM_isZero ? 28'h0 : _T_678; // @[Mux.scala 87:16]
  assign io_M = decM_isNaR ? 28'h8000000 : _T_680; // @[PositMultiplier.scala 86:8]
endmodule
