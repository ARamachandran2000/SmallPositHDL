module PositFMA28_3(
  input         clock,
  input         reset,
  input         io_inValid,
  input  [1:0]  io_fmaOp,
  input  [27:0] io_A,
  input  [27:0] io_B,
  input  [27:0] io_C,
  output [27:0] io_F,
  output        io_outValid
);
  wire  _T; // @[PositFMA.scala 47:36]
  wire [27:0] _T_2; // @[Bitwise.scala 71:12]
  wire [27:0] _T_3; // @[PositFMA.scala 47:41]
  wire [27:0] _GEN_10; // @[PositFMA.scala 47:49]
  wire [27:0] realA; // @[PositFMA.scala 47:49]
  wire  _T_6; // @[PositFMA.scala 48:36]
  wire [27:0] _T_8; // @[Bitwise.scala 71:12]
  wire [27:0] _T_9; // @[PositFMA.scala 48:41]
  wire [27:0] _GEN_11; // @[PositFMA.scala 48:49]
  wire [27:0] realC; // @[PositFMA.scala 48:49]
  wire  _T_13; // @[convert.scala 18:24]
  wire  _T_14; // @[convert.scala 18:40]
  wire  _T_15; // @[convert.scala 18:36]
  wire [25:0] _T_16; // @[convert.scala 19:24]
  wire [25:0] _T_17; // @[convert.scala 19:43]
  wire [25:0] _T_18; // @[convert.scala 19:39]
  wire [15:0] _T_19; // @[LZD.scala 43:32]
  wire [7:0] _T_20; // @[LZD.scala 43:32]
  wire [3:0] _T_21; // @[LZD.scala 43:32]
  wire [1:0] _T_22; // @[LZD.scala 43:32]
  wire  _T_23; // @[LZD.scala 39:14]
  wire  _T_24; // @[LZD.scala 39:21]
  wire  _T_25; // @[LZD.scala 39:30]
  wire  _T_26; // @[LZD.scala 39:27]
  wire  _T_27; // @[LZD.scala 39:25]
  wire [1:0] _T_28; // @[Cat.scala 29:58]
  wire [1:0] _T_29; // @[LZD.scala 44:32]
  wire  _T_30; // @[LZD.scala 39:14]
  wire  _T_31; // @[LZD.scala 39:21]
  wire  _T_32; // @[LZD.scala 39:30]
  wire  _T_33; // @[LZD.scala 39:27]
  wire  _T_34; // @[LZD.scala 39:25]
  wire [1:0] _T_35; // @[Cat.scala 29:58]
  wire  _T_36; // @[Shift.scala 12:21]
  wire  _T_37; // @[Shift.scala 12:21]
  wire  _T_38; // @[LZD.scala 49:16]
  wire  _T_39; // @[LZD.scala 49:27]
  wire  _T_40; // @[LZD.scala 49:25]
  wire  _T_41; // @[LZD.scala 49:47]
  wire  _T_42; // @[LZD.scala 49:59]
  wire  _T_43; // @[LZD.scala 49:35]
  wire [2:0] _T_45; // @[Cat.scala 29:58]
  wire [3:0] _T_46; // @[LZD.scala 44:32]
  wire [1:0] _T_47; // @[LZD.scala 43:32]
  wire  _T_48; // @[LZD.scala 39:14]
  wire  _T_49; // @[LZD.scala 39:21]
  wire  _T_50; // @[LZD.scala 39:30]
  wire  _T_51; // @[LZD.scala 39:27]
  wire  _T_52; // @[LZD.scala 39:25]
  wire [1:0] _T_53; // @[Cat.scala 29:58]
  wire [1:0] _T_54; // @[LZD.scala 44:32]
  wire  _T_55; // @[LZD.scala 39:14]
  wire  _T_56; // @[LZD.scala 39:21]
  wire  _T_57; // @[LZD.scala 39:30]
  wire  _T_58; // @[LZD.scala 39:27]
  wire  _T_59; // @[LZD.scala 39:25]
  wire [1:0] _T_60; // @[Cat.scala 29:58]
  wire  _T_61; // @[Shift.scala 12:21]
  wire  _T_62; // @[Shift.scala 12:21]
  wire  _T_63; // @[LZD.scala 49:16]
  wire  _T_64; // @[LZD.scala 49:27]
  wire  _T_65; // @[LZD.scala 49:25]
  wire  _T_66; // @[LZD.scala 49:47]
  wire  _T_67; // @[LZD.scala 49:59]
  wire  _T_68; // @[LZD.scala 49:35]
  wire [2:0] _T_70; // @[Cat.scala 29:58]
  wire  _T_71; // @[Shift.scala 12:21]
  wire  _T_72; // @[Shift.scala 12:21]
  wire  _T_73; // @[LZD.scala 49:16]
  wire  _T_74; // @[LZD.scala 49:27]
  wire  _T_75; // @[LZD.scala 49:25]
  wire [1:0] _T_76; // @[LZD.scala 49:47]
  wire [1:0] _T_77; // @[LZD.scala 49:59]
  wire [1:0] _T_78; // @[LZD.scala 49:35]
  wire [3:0] _T_80; // @[Cat.scala 29:58]
  wire [7:0] _T_81; // @[LZD.scala 44:32]
  wire [3:0] _T_82; // @[LZD.scala 43:32]
  wire [1:0] _T_83; // @[LZD.scala 43:32]
  wire  _T_84; // @[LZD.scala 39:14]
  wire  _T_85; // @[LZD.scala 39:21]
  wire  _T_86; // @[LZD.scala 39:30]
  wire  _T_87; // @[LZD.scala 39:27]
  wire  _T_88; // @[LZD.scala 39:25]
  wire [1:0] _T_89; // @[Cat.scala 29:58]
  wire [1:0] _T_90; // @[LZD.scala 44:32]
  wire  _T_91; // @[LZD.scala 39:14]
  wire  _T_92; // @[LZD.scala 39:21]
  wire  _T_93; // @[LZD.scala 39:30]
  wire  _T_94; // @[LZD.scala 39:27]
  wire  _T_95; // @[LZD.scala 39:25]
  wire [1:0] _T_96; // @[Cat.scala 29:58]
  wire  _T_97; // @[Shift.scala 12:21]
  wire  _T_98; // @[Shift.scala 12:21]
  wire  _T_99; // @[LZD.scala 49:16]
  wire  _T_100; // @[LZD.scala 49:27]
  wire  _T_101; // @[LZD.scala 49:25]
  wire  _T_102; // @[LZD.scala 49:47]
  wire  _T_103; // @[LZD.scala 49:59]
  wire  _T_104; // @[LZD.scala 49:35]
  wire [2:0] _T_106; // @[Cat.scala 29:58]
  wire [3:0] _T_107; // @[LZD.scala 44:32]
  wire [1:0] _T_108; // @[LZD.scala 43:32]
  wire  _T_109; // @[LZD.scala 39:14]
  wire  _T_110; // @[LZD.scala 39:21]
  wire  _T_111; // @[LZD.scala 39:30]
  wire  _T_112; // @[LZD.scala 39:27]
  wire  _T_113; // @[LZD.scala 39:25]
  wire [1:0] _T_114; // @[Cat.scala 29:58]
  wire [1:0] _T_115; // @[LZD.scala 44:32]
  wire  _T_116; // @[LZD.scala 39:14]
  wire  _T_117; // @[LZD.scala 39:21]
  wire  _T_118; // @[LZD.scala 39:30]
  wire  _T_119; // @[LZD.scala 39:27]
  wire  _T_120; // @[LZD.scala 39:25]
  wire [1:0] _T_121; // @[Cat.scala 29:58]
  wire  _T_122; // @[Shift.scala 12:21]
  wire  _T_123; // @[Shift.scala 12:21]
  wire  _T_124; // @[LZD.scala 49:16]
  wire  _T_125; // @[LZD.scala 49:27]
  wire  _T_126; // @[LZD.scala 49:25]
  wire  _T_127; // @[LZD.scala 49:47]
  wire  _T_128; // @[LZD.scala 49:59]
  wire  _T_129; // @[LZD.scala 49:35]
  wire [2:0] _T_131; // @[Cat.scala 29:58]
  wire  _T_132; // @[Shift.scala 12:21]
  wire  _T_133; // @[Shift.scala 12:21]
  wire  _T_134; // @[LZD.scala 49:16]
  wire  _T_135; // @[LZD.scala 49:27]
  wire  _T_136; // @[LZD.scala 49:25]
  wire [1:0] _T_137; // @[LZD.scala 49:47]
  wire [1:0] _T_138; // @[LZD.scala 49:59]
  wire [1:0] _T_139; // @[LZD.scala 49:35]
  wire [3:0] _T_141; // @[Cat.scala 29:58]
  wire  _T_142; // @[Shift.scala 12:21]
  wire  _T_143; // @[Shift.scala 12:21]
  wire  _T_144; // @[LZD.scala 49:16]
  wire  _T_145; // @[LZD.scala 49:27]
  wire  _T_146; // @[LZD.scala 49:25]
  wire [2:0] _T_147; // @[LZD.scala 49:47]
  wire [2:0] _T_148; // @[LZD.scala 49:59]
  wire [2:0] _T_149; // @[LZD.scala 49:35]
  wire [4:0] _T_151; // @[Cat.scala 29:58]
  wire [9:0] _T_152; // @[LZD.scala 44:32]
  wire [7:0] _T_153; // @[LZD.scala 43:32]
  wire [3:0] _T_154; // @[LZD.scala 43:32]
  wire [1:0] _T_155; // @[LZD.scala 43:32]
  wire  _T_156; // @[LZD.scala 39:14]
  wire  _T_157; // @[LZD.scala 39:21]
  wire  _T_158; // @[LZD.scala 39:30]
  wire  _T_159; // @[LZD.scala 39:27]
  wire  _T_160; // @[LZD.scala 39:25]
  wire [1:0] _T_161; // @[Cat.scala 29:58]
  wire [1:0] _T_162; // @[LZD.scala 44:32]
  wire  _T_163; // @[LZD.scala 39:14]
  wire  _T_164; // @[LZD.scala 39:21]
  wire  _T_165; // @[LZD.scala 39:30]
  wire  _T_166; // @[LZD.scala 39:27]
  wire  _T_167; // @[LZD.scala 39:25]
  wire [1:0] _T_168; // @[Cat.scala 29:58]
  wire  _T_169; // @[Shift.scala 12:21]
  wire  _T_170; // @[Shift.scala 12:21]
  wire  _T_171; // @[LZD.scala 49:16]
  wire  _T_172; // @[LZD.scala 49:27]
  wire  _T_173; // @[LZD.scala 49:25]
  wire  _T_174; // @[LZD.scala 49:47]
  wire  _T_175; // @[LZD.scala 49:59]
  wire  _T_176; // @[LZD.scala 49:35]
  wire [2:0] _T_178; // @[Cat.scala 29:58]
  wire [3:0] _T_179; // @[LZD.scala 44:32]
  wire [1:0] _T_180; // @[LZD.scala 43:32]
  wire  _T_181; // @[LZD.scala 39:14]
  wire  _T_182; // @[LZD.scala 39:21]
  wire  _T_183; // @[LZD.scala 39:30]
  wire  _T_184; // @[LZD.scala 39:27]
  wire  _T_185; // @[LZD.scala 39:25]
  wire [1:0] _T_186; // @[Cat.scala 29:58]
  wire [1:0] _T_187; // @[LZD.scala 44:32]
  wire  _T_188; // @[LZD.scala 39:14]
  wire  _T_189; // @[LZD.scala 39:21]
  wire  _T_190; // @[LZD.scala 39:30]
  wire  _T_191; // @[LZD.scala 39:27]
  wire  _T_192; // @[LZD.scala 39:25]
  wire [1:0] _T_193; // @[Cat.scala 29:58]
  wire  _T_194; // @[Shift.scala 12:21]
  wire  _T_195; // @[Shift.scala 12:21]
  wire  _T_196; // @[LZD.scala 49:16]
  wire  _T_197; // @[LZD.scala 49:27]
  wire  _T_198; // @[LZD.scala 49:25]
  wire  _T_199; // @[LZD.scala 49:47]
  wire  _T_200; // @[LZD.scala 49:59]
  wire  _T_201; // @[LZD.scala 49:35]
  wire [2:0] _T_203; // @[Cat.scala 29:58]
  wire  _T_204; // @[Shift.scala 12:21]
  wire  _T_205; // @[Shift.scala 12:21]
  wire  _T_206; // @[LZD.scala 49:16]
  wire  _T_207; // @[LZD.scala 49:27]
  wire  _T_208; // @[LZD.scala 49:25]
  wire [1:0] _T_209; // @[LZD.scala 49:47]
  wire [1:0] _T_210; // @[LZD.scala 49:59]
  wire [1:0] _T_211; // @[LZD.scala 49:35]
  wire [3:0] _T_213; // @[Cat.scala 29:58]
  wire [1:0] _T_214; // @[LZD.scala 44:32]
  wire  _T_215; // @[LZD.scala 39:14]
  wire  _T_216; // @[LZD.scala 39:21]
  wire  _T_217; // @[LZD.scala 39:30]
  wire  _T_218; // @[LZD.scala 39:27]
  wire  _T_219; // @[LZD.scala 39:25]
  wire  _T_221; // @[Shift.scala 12:21]
  wire [2:0] _T_223; // @[Cat.scala 29:58]
  wire [2:0] _T_224; // @[LZD.scala 55:32]
  wire [2:0] _T_225; // @[LZD.scala 55:20]
  wire [3:0] _T_226; // @[Cat.scala 29:58]
  wire  _T_227; // @[Shift.scala 12:21]
  wire [3:0] _T_229; // @[LZD.scala 55:32]
  wire [3:0] _T_230; // @[LZD.scala 55:20]
  wire [4:0] _T_231; // @[Cat.scala 29:58]
  wire [4:0] _T_232; // @[convert.scala 21:22]
  wire [24:0] _T_233; // @[convert.scala 22:36]
  wire  _T_234; // @[Shift.scala 16:24]
  wire  _T_236; // @[Shift.scala 12:21]
  wire [8:0] _T_237; // @[Shift.scala 64:52]
  wire [24:0] _T_239; // @[Cat.scala 29:58]
  wire [24:0] _T_240; // @[Shift.scala 64:27]
  wire [3:0] _T_241; // @[Shift.scala 66:70]
  wire  _T_242; // @[Shift.scala 12:21]
  wire [16:0] _T_243; // @[Shift.scala 64:52]
  wire [24:0] _T_245; // @[Cat.scala 29:58]
  wire [24:0] _T_246; // @[Shift.scala 64:27]
  wire [2:0] _T_247; // @[Shift.scala 66:70]
  wire  _T_248; // @[Shift.scala 12:21]
  wire [20:0] _T_249; // @[Shift.scala 64:52]
  wire [24:0] _T_251; // @[Cat.scala 29:58]
  wire [24:0] _T_252; // @[Shift.scala 64:27]
  wire [1:0] _T_253; // @[Shift.scala 66:70]
  wire  _T_254; // @[Shift.scala 12:21]
  wire [22:0] _T_255; // @[Shift.scala 64:52]
  wire [24:0] _T_257; // @[Cat.scala 29:58]
  wire [24:0] _T_258; // @[Shift.scala 64:27]
  wire  _T_259; // @[Shift.scala 66:70]
  wire [23:0] _T_261; // @[Shift.scala 64:52]
  wire [24:0] _T_262; // @[Cat.scala 29:58]
  wire [24:0] _T_263; // @[Shift.scala 64:27]
  wire [24:0] _T_264; // @[Shift.scala 16:10]
  wire [2:0] _T_265; // @[convert.scala 23:34]
  wire [21:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_267; // @[convert.scala 25:26]
  wire [4:0] _T_269; // @[convert.scala 25:42]
  wire [2:0] _T_272; // @[convert.scala 26:67]
  wire [2:0] _T_273; // @[convert.scala 26:51]
  wire [8:0] _T_274; // @[Cat.scala 29:58]
  wire [26:0] _T_276; // @[convert.scala 29:56]
  wire  _T_277; // @[convert.scala 29:60]
  wire  _T_278; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_281; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [8:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_290; // @[convert.scala 18:24]
  wire  _T_291; // @[convert.scala 18:40]
  wire  _T_292; // @[convert.scala 18:36]
  wire [25:0] _T_293; // @[convert.scala 19:24]
  wire [25:0] _T_294; // @[convert.scala 19:43]
  wire [25:0] _T_295; // @[convert.scala 19:39]
  wire [15:0] _T_296; // @[LZD.scala 43:32]
  wire [7:0] _T_297; // @[LZD.scala 43:32]
  wire [3:0] _T_298; // @[LZD.scala 43:32]
  wire [1:0] _T_299; // @[LZD.scala 43:32]
  wire  _T_300; // @[LZD.scala 39:14]
  wire  _T_301; // @[LZD.scala 39:21]
  wire  _T_302; // @[LZD.scala 39:30]
  wire  _T_303; // @[LZD.scala 39:27]
  wire  _T_304; // @[LZD.scala 39:25]
  wire [1:0] _T_305; // @[Cat.scala 29:58]
  wire [1:0] _T_306; // @[LZD.scala 44:32]
  wire  _T_307; // @[LZD.scala 39:14]
  wire  _T_308; // @[LZD.scala 39:21]
  wire  _T_309; // @[LZD.scala 39:30]
  wire  _T_310; // @[LZD.scala 39:27]
  wire  _T_311; // @[LZD.scala 39:25]
  wire [1:0] _T_312; // @[Cat.scala 29:58]
  wire  _T_313; // @[Shift.scala 12:21]
  wire  _T_314; // @[Shift.scala 12:21]
  wire  _T_315; // @[LZD.scala 49:16]
  wire  _T_316; // @[LZD.scala 49:27]
  wire  _T_317; // @[LZD.scala 49:25]
  wire  _T_318; // @[LZD.scala 49:47]
  wire  _T_319; // @[LZD.scala 49:59]
  wire  _T_320; // @[LZD.scala 49:35]
  wire [2:0] _T_322; // @[Cat.scala 29:58]
  wire [3:0] _T_323; // @[LZD.scala 44:32]
  wire [1:0] _T_324; // @[LZD.scala 43:32]
  wire  _T_325; // @[LZD.scala 39:14]
  wire  _T_326; // @[LZD.scala 39:21]
  wire  _T_327; // @[LZD.scala 39:30]
  wire  _T_328; // @[LZD.scala 39:27]
  wire  _T_329; // @[LZD.scala 39:25]
  wire [1:0] _T_330; // @[Cat.scala 29:58]
  wire [1:0] _T_331; // @[LZD.scala 44:32]
  wire  _T_332; // @[LZD.scala 39:14]
  wire  _T_333; // @[LZD.scala 39:21]
  wire  _T_334; // @[LZD.scala 39:30]
  wire  _T_335; // @[LZD.scala 39:27]
  wire  _T_336; // @[LZD.scala 39:25]
  wire [1:0] _T_337; // @[Cat.scala 29:58]
  wire  _T_338; // @[Shift.scala 12:21]
  wire  _T_339; // @[Shift.scala 12:21]
  wire  _T_340; // @[LZD.scala 49:16]
  wire  _T_341; // @[LZD.scala 49:27]
  wire  _T_342; // @[LZD.scala 49:25]
  wire  _T_343; // @[LZD.scala 49:47]
  wire  _T_344; // @[LZD.scala 49:59]
  wire  _T_345; // @[LZD.scala 49:35]
  wire [2:0] _T_347; // @[Cat.scala 29:58]
  wire  _T_348; // @[Shift.scala 12:21]
  wire  _T_349; // @[Shift.scala 12:21]
  wire  _T_350; // @[LZD.scala 49:16]
  wire  _T_351; // @[LZD.scala 49:27]
  wire  _T_352; // @[LZD.scala 49:25]
  wire [1:0] _T_353; // @[LZD.scala 49:47]
  wire [1:0] _T_354; // @[LZD.scala 49:59]
  wire [1:0] _T_355; // @[LZD.scala 49:35]
  wire [3:0] _T_357; // @[Cat.scala 29:58]
  wire [7:0] _T_358; // @[LZD.scala 44:32]
  wire [3:0] _T_359; // @[LZD.scala 43:32]
  wire [1:0] _T_360; // @[LZD.scala 43:32]
  wire  _T_361; // @[LZD.scala 39:14]
  wire  _T_362; // @[LZD.scala 39:21]
  wire  _T_363; // @[LZD.scala 39:30]
  wire  _T_364; // @[LZD.scala 39:27]
  wire  _T_365; // @[LZD.scala 39:25]
  wire [1:0] _T_366; // @[Cat.scala 29:58]
  wire [1:0] _T_367; // @[LZD.scala 44:32]
  wire  _T_368; // @[LZD.scala 39:14]
  wire  _T_369; // @[LZD.scala 39:21]
  wire  _T_370; // @[LZD.scala 39:30]
  wire  _T_371; // @[LZD.scala 39:27]
  wire  _T_372; // @[LZD.scala 39:25]
  wire [1:0] _T_373; // @[Cat.scala 29:58]
  wire  _T_374; // @[Shift.scala 12:21]
  wire  _T_375; // @[Shift.scala 12:21]
  wire  _T_376; // @[LZD.scala 49:16]
  wire  _T_377; // @[LZD.scala 49:27]
  wire  _T_378; // @[LZD.scala 49:25]
  wire  _T_379; // @[LZD.scala 49:47]
  wire  _T_380; // @[LZD.scala 49:59]
  wire  _T_381; // @[LZD.scala 49:35]
  wire [2:0] _T_383; // @[Cat.scala 29:58]
  wire [3:0] _T_384; // @[LZD.scala 44:32]
  wire [1:0] _T_385; // @[LZD.scala 43:32]
  wire  _T_386; // @[LZD.scala 39:14]
  wire  _T_387; // @[LZD.scala 39:21]
  wire  _T_388; // @[LZD.scala 39:30]
  wire  _T_389; // @[LZD.scala 39:27]
  wire  _T_390; // @[LZD.scala 39:25]
  wire [1:0] _T_391; // @[Cat.scala 29:58]
  wire [1:0] _T_392; // @[LZD.scala 44:32]
  wire  _T_393; // @[LZD.scala 39:14]
  wire  _T_394; // @[LZD.scala 39:21]
  wire  _T_395; // @[LZD.scala 39:30]
  wire  _T_396; // @[LZD.scala 39:27]
  wire  _T_397; // @[LZD.scala 39:25]
  wire [1:0] _T_398; // @[Cat.scala 29:58]
  wire  _T_399; // @[Shift.scala 12:21]
  wire  _T_400; // @[Shift.scala 12:21]
  wire  _T_401; // @[LZD.scala 49:16]
  wire  _T_402; // @[LZD.scala 49:27]
  wire  _T_403; // @[LZD.scala 49:25]
  wire  _T_404; // @[LZD.scala 49:47]
  wire  _T_405; // @[LZD.scala 49:59]
  wire  _T_406; // @[LZD.scala 49:35]
  wire [2:0] _T_408; // @[Cat.scala 29:58]
  wire  _T_409; // @[Shift.scala 12:21]
  wire  _T_410; // @[Shift.scala 12:21]
  wire  _T_411; // @[LZD.scala 49:16]
  wire  _T_412; // @[LZD.scala 49:27]
  wire  _T_413; // @[LZD.scala 49:25]
  wire [1:0] _T_414; // @[LZD.scala 49:47]
  wire [1:0] _T_415; // @[LZD.scala 49:59]
  wire [1:0] _T_416; // @[LZD.scala 49:35]
  wire [3:0] _T_418; // @[Cat.scala 29:58]
  wire  _T_419; // @[Shift.scala 12:21]
  wire  _T_420; // @[Shift.scala 12:21]
  wire  _T_421; // @[LZD.scala 49:16]
  wire  _T_422; // @[LZD.scala 49:27]
  wire  _T_423; // @[LZD.scala 49:25]
  wire [2:0] _T_424; // @[LZD.scala 49:47]
  wire [2:0] _T_425; // @[LZD.scala 49:59]
  wire [2:0] _T_426; // @[LZD.scala 49:35]
  wire [4:0] _T_428; // @[Cat.scala 29:58]
  wire [9:0] _T_429; // @[LZD.scala 44:32]
  wire [7:0] _T_430; // @[LZD.scala 43:32]
  wire [3:0] _T_431; // @[LZD.scala 43:32]
  wire [1:0] _T_432; // @[LZD.scala 43:32]
  wire  _T_433; // @[LZD.scala 39:14]
  wire  _T_434; // @[LZD.scala 39:21]
  wire  _T_435; // @[LZD.scala 39:30]
  wire  _T_436; // @[LZD.scala 39:27]
  wire  _T_437; // @[LZD.scala 39:25]
  wire [1:0] _T_438; // @[Cat.scala 29:58]
  wire [1:0] _T_439; // @[LZD.scala 44:32]
  wire  _T_440; // @[LZD.scala 39:14]
  wire  _T_441; // @[LZD.scala 39:21]
  wire  _T_442; // @[LZD.scala 39:30]
  wire  _T_443; // @[LZD.scala 39:27]
  wire  _T_444; // @[LZD.scala 39:25]
  wire [1:0] _T_445; // @[Cat.scala 29:58]
  wire  _T_446; // @[Shift.scala 12:21]
  wire  _T_447; // @[Shift.scala 12:21]
  wire  _T_448; // @[LZD.scala 49:16]
  wire  _T_449; // @[LZD.scala 49:27]
  wire  _T_450; // @[LZD.scala 49:25]
  wire  _T_451; // @[LZD.scala 49:47]
  wire  _T_452; // @[LZD.scala 49:59]
  wire  _T_453; // @[LZD.scala 49:35]
  wire [2:0] _T_455; // @[Cat.scala 29:58]
  wire [3:0] _T_456; // @[LZD.scala 44:32]
  wire [1:0] _T_457; // @[LZD.scala 43:32]
  wire  _T_458; // @[LZD.scala 39:14]
  wire  _T_459; // @[LZD.scala 39:21]
  wire  _T_460; // @[LZD.scala 39:30]
  wire  _T_461; // @[LZD.scala 39:27]
  wire  _T_462; // @[LZD.scala 39:25]
  wire [1:0] _T_463; // @[Cat.scala 29:58]
  wire [1:0] _T_464; // @[LZD.scala 44:32]
  wire  _T_465; // @[LZD.scala 39:14]
  wire  _T_466; // @[LZD.scala 39:21]
  wire  _T_467; // @[LZD.scala 39:30]
  wire  _T_468; // @[LZD.scala 39:27]
  wire  _T_469; // @[LZD.scala 39:25]
  wire [1:0] _T_470; // @[Cat.scala 29:58]
  wire  _T_471; // @[Shift.scala 12:21]
  wire  _T_472; // @[Shift.scala 12:21]
  wire  _T_473; // @[LZD.scala 49:16]
  wire  _T_474; // @[LZD.scala 49:27]
  wire  _T_475; // @[LZD.scala 49:25]
  wire  _T_476; // @[LZD.scala 49:47]
  wire  _T_477; // @[LZD.scala 49:59]
  wire  _T_478; // @[LZD.scala 49:35]
  wire [2:0] _T_480; // @[Cat.scala 29:58]
  wire  _T_481; // @[Shift.scala 12:21]
  wire  _T_482; // @[Shift.scala 12:21]
  wire  _T_483; // @[LZD.scala 49:16]
  wire  _T_484; // @[LZD.scala 49:27]
  wire  _T_485; // @[LZD.scala 49:25]
  wire [1:0] _T_486; // @[LZD.scala 49:47]
  wire [1:0] _T_487; // @[LZD.scala 49:59]
  wire [1:0] _T_488; // @[LZD.scala 49:35]
  wire [3:0] _T_490; // @[Cat.scala 29:58]
  wire [1:0] _T_491; // @[LZD.scala 44:32]
  wire  _T_492; // @[LZD.scala 39:14]
  wire  _T_493; // @[LZD.scala 39:21]
  wire  _T_494; // @[LZD.scala 39:30]
  wire  _T_495; // @[LZD.scala 39:27]
  wire  _T_496; // @[LZD.scala 39:25]
  wire  _T_498; // @[Shift.scala 12:21]
  wire [2:0] _T_500; // @[Cat.scala 29:58]
  wire [2:0] _T_501; // @[LZD.scala 55:32]
  wire [2:0] _T_502; // @[LZD.scala 55:20]
  wire [3:0] _T_503; // @[Cat.scala 29:58]
  wire  _T_504; // @[Shift.scala 12:21]
  wire [3:0] _T_506; // @[LZD.scala 55:32]
  wire [3:0] _T_507; // @[LZD.scala 55:20]
  wire [4:0] _T_508; // @[Cat.scala 29:58]
  wire [4:0] _T_509; // @[convert.scala 21:22]
  wire [24:0] _T_510; // @[convert.scala 22:36]
  wire  _T_511; // @[Shift.scala 16:24]
  wire  _T_513; // @[Shift.scala 12:21]
  wire [8:0] _T_514; // @[Shift.scala 64:52]
  wire [24:0] _T_516; // @[Cat.scala 29:58]
  wire [24:0] _T_517; // @[Shift.scala 64:27]
  wire [3:0] _T_518; // @[Shift.scala 66:70]
  wire  _T_519; // @[Shift.scala 12:21]
  wire [16:0] _T_520; // @[Shift.scala 64:52]
  wire [24:0] _T_522; // @[Cat.scala 29:58]
  wire [24:0] _T_523; // @[Shift.scala 64:27]
  wire [2:0] _T_524; // @[Shift.scala 66:70]
  wire  _T_525; // @[Shift.scala 12:21]
  wire [20:0] _T_526; // @[Shift.scala 64:52]
  wire [24:0] _T_528; // @[Cat.scala 29:58]
  wire [24:0] _T_529; // @[Shift.scala 64:27]
  wire [1:0] _T_530; // @[Shift.scala 66:70]
  wire  _T_531; // @[Shift.scala 12:21]
  wire [22:0] _T_532; // @[Shift.scala 64:52]
  wire [24:0] _T_534; // @[Cat.scala 29:58]
  wire [24:0] _T_535; // @[Shift.scala 64:27]
  wire  _T_536; // @[Shift.scala 66:70]
  wire [23:0] _T_538; // @[Shift.scala 64:52]
  wire [24:0] _T_539; // @[Cat.scala 29:58]
  wire [24:0] _T_540; // @[Shift.scala 64:27]
  wire [24:0] _T_541; // @[Shift.scala 16:10]
  wire [2:0] _T_542; // @[convert.scala 23:34]
  wire [21:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_544; // @[convert.scala 25:26]
  wire [4:0] _T_546; // @[convert.scala 25:42]
  wire [2:0] _T_549; // @[convert.scala 26:67]
  wire [2:0] _T_550; // @[convert.scala 26:51]
  wire [8:0] _T_551; // @[Cat.scala 29:58]
  wire [26:0] _T_553; // @[convert.scala 29:56]
  wire  _T_554; // @[convert.scala 29:60]
  wire  _T_555; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_558; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [8:0] decB_scale; // @[convert.scala 32:24]
  wire  _T_567; // @[convert.scala 18:24]
  wire  _T_568; // @[convert.scala 18:40]
  wire  _T_569; // @[convert.scala 18:36]
  wire [25:0] _T_570; // @[convert.scala 19:24]
  wire [25:0] _T_571; // @[convert.scala 19:43]
  wire [25:0] _T_572; // @[convert.scala 19:39]
  wire [15:0] _T_573; // @[LZD.scala 43:32]
  wire [7:0] _T_574; // @[LZD.scala 43:32]
  wire [3:0] _T_575; // @[LZD.scala 43:32]
  wire [1:0] _T_576; // @[LZD.scala 43:32]
  wire  _T_577; // @[LZD.scala 39:14]
  wire  _T_578; // @[LZD.scala 39:21]
  wire  _T_579; // @[LZD.scala 39:30]
  wire  _T_580; // @[LZD.scala 39:27]
  wire  _T_581; // @[LZD.scala 39:25]
  wire [1:0] _T_582; // @[Cat.scala 29:58]
  wire [1:0] _T_583; // @[LZD.scala 44:32]
  wire  _T_584; // @[LZD.scala 39:14]
  wire  _T_585; // @[LZD.scala 39:21]
  wire  _T_586; // @[LZD.scala 39:30]
  wire  _T_587; // @[LZD.scala 39:27]
  wire  _T_588; // @[LZD.scala 39:25]
  wire [1:0] _T_589; // @[Cat.scala 29:58]
  wire  _T_590; // @[Shift.scala 12:21]
  wire  _T_591; // @[Shift.scala 12:21]
  wire  _T_592; // @[LZD.scala 49:16]
  wire  _T_593; // @[LZD.scala 49:27]
  wire  _T_594; // @[LZD.scala 49:25]
  wire  _T_595; // @[LZD.scala 49:47]
  wire  _T_596; // @[LZD.scala 49:59]
  wire  _T_597; // @[LZD.scala 49:35]
  wire [2:0] _T_599; // @[Cat.scala 29:58]
  wire [3:0] _T_600; // @[LZD.scala 44:32]
  wire [1:0] _T_601; // @[LZD.scala 43:32]
  wire  _T_602; // @[LZD.scala 39:14]
  wire  _T_603; // @[LZD.scala 39:21]
  wire  _T_604; // @[LZD.scala 39:30]
  wire  _T_605; // @[LZD.scala 39:27]
  wire  _T_606; // @[LZD.scala 39:25]
  wire [1:0] _T_607; // @[Cat.scala 29:58]
  wire [1:0] _T_608; // @[LZD.scala 44:32]
  wire  _T_609; // @[LZD.scala 39:14]
  wire  _T_610; // @[LZD.scala 39:21]
  wire  _T_611; // @[LZD.scala 39:30]
  wire  _T_612; // @[LZD.scala 39:27]
  wire  _T_613; // @[LZD.scala 39:25]
  wire [1:0] _T_614; // @[Cat.scala 29:58]
  wire  _T_615; // @[Shift.scala 12:21]
  wire  _T_616; // @[Shift.scala 12:21]
  wire  _T_617; // @[LZD.scala 49:16]
  wire  _T_618; // @[LZD.scala 49:27]
  wire  _T_619; // @[LZD.scala 49:25]
  wire  _T_620; // @[LZD.scala 49:47]
  wire  _T_621; // @[LZD.scala 49:59]
  wire  _T_622; // @[LZD.scala 49:35]
  wire [2:0] _T_624; // @[Cat.scala 29:58]
  wire  _T_625; // @[Shift.scala 12:21]
  wire  _T_626; // @[Shift.scala 12:21]
  wire  _T_627; // @[LZD.scala 49:16]
  wire  _T_628; // @[LZD.scala 49:27]
  wire  _T_629; // @[LZD.scala 49:25]
  wire [1:0] _T_630; // @[LZD.scala 49:47]
  wire [1:0] _T_631; // @[LZD.scala 49:59]
  wire [1:0] _T_632; // @[LZD.scala 49:35]
  wire [3:0] _T_634; // @[Cat.scala 29:58]
  wire [7:0] _T_635; // @[LZD.scala 44:32]
  wire [3:0] _T_636; // @[LZD.scala 43:32]
  wire [1:0] _T_637; // @[LZD.scala 43:32]
  wire  _T_638; // @[LZD.scala 39:14]
  wire  _T_639; // @[LZD.scala 39:21]
  wire  _T_640; // @[LZD.scala 39:30]
  wire  _T_641; // @[LZD.scala 39:27]
  wire  _T_642; // @[LZD.scala 39:25]
  wire [1:0] _T_643; // @[Cat.scala 29:58]
  wire [1:0] _T_644; // @[LZD.scala 44:32]
  wire  _T_645; // @[LZD.scala 39:14]
  wire  _T_646; // @[LZD.scala 39:21]
  wire  _T_647; // @[LZD.scala 39:30]
  wire  _T_648; // @[LZD.scala 39:27]
  wire  _T_649; // @[LZD.scala 39:25]
  wire [1:0] _T_650; // @[Cat.scala 29:58]
  wire  _T_651; // @[Shift.scala 12:21]
  wire  _T_652; // @[Shift.scala 12:21]
  wire  _T_653; // @[LZD.scala 49:16]
  wire  _T_654; // @[LZD.scala 49:27]
  wire  _T_655; // @[LZD.scala 49:25]
  wire  _T_656; // @[LZD.scala 49:47]
  wire  _T_657; // @[LZD.scala 49:59]
  wire  _T_658; // @[LZD.scala 49:35]
  wire [2:0] _T_660; // @[Cat.scala 29:58]
  wire [3:0] _T_661; // @[LZD.scala 44:32]
  wire [1:0] _T_662; // @[LZD.scala 43:32]
  wire  _T_663; // @[LZD.scala 39:14]
  wire  _T_664; // @[LZD.scala 39:21]
  wire  _T_665; // @[LZD.scala 39:30]
  wire  _T_666; // @[LZD.scala 39:27]
  wire  _T_667; // @[LZD.scala 39:25]
  wire [1:0] _T_668; // @[Cat.scala 29:58]
  wire [1:0] _T_669; // @[LZD.scala 44:32]
  wire  _T_670; // @[LZD.scala 39:14]
  wire  _T_671; // @[LZD.scala 39:21]
  wire  _T_672; // @[LZD.scala 39:30]
  wire  _T_673; // @[LZD.scala 39:27]
  wire  _T_674; // @[LZD.scala 39:25]
  wire [1:0] _T_675; // @[Cat.scala 29:58]
  wire  _T_676; // @[Shift.scala 12:21]
  wire  _T_677; // @[Shift.scala 12:21]
  wire  _T_678; // @[LZD.scala 49:16]
  wire  _T_679; // @[LZD.scala 49:27]
  wire  _T_680; // @[LZD.scala 49:25]
  wire  _T_681; // @[LZD.scala 49:47]
  wire  _T_682; // @[LZD.scala 49:59]
  wire  _T_683; // @[LZD.scala 49:35]
  wire [2:0] _T_685; // @[Cat.scala 29:58]
  wire  _T_686; // @[Shift.scala 12:21]
  wire  _T_687; // @[Shift.scala 12:21]
  wire  _T_688; // @[LZD.scala 49:16]
  wire  _T_689; // @[LZD.scala 49:27]
  wire  _T_690; // @[LZD.scala 49:25]
  wire [1:0] _T_691; // @[LZD.scala 49:47]
  wire [1:0] _T_692; // @[LZD.scala 49:59]
  wire [1:0] _T_693; // @[LZD.scala 49:35]
  wire [3:0] _T_695; // @[Cat.scala 29:58]
  wire  _T_696; // @[Shift.scala 12:21]
  wire  _T_697; // @[Shift.scala 12:21]
  wire  _T_698; // @[LZD.scala 49:16]
  wire  _T_699; // @[LZD.scala 49:27]
  wire  _T_700; // @[LZD.scala 49:25]
  wire [2:0] _T_701; // @[LZD.scala 49:47]
  wire [2:0] _T_702; // @[LZD.scala 49:59]
  wire [2:0] _T_703; // @[LZD.scala 49:35]
  wire [4:0] _T_705; // @[Cat.scala 29:58]
  wire [9:0] _T_706; // @[LZD.scala 44:32]
  wire [7:0] _T_707; // @[LZD.scala 43:32]
  wire [3:0] _T_708; // @[LZD.scala 43:32]
  wire [1:0] _T_709; // @[LZD.scala 43:32]
  wire  _T_710; // @[LZD.scala 39:14]
  wire  _T_711; // @[LZD.scala 39:21]
  wire  _T_712; // @[LZD.scala 39:30]
  wire  _T_713; // @[LZD.scala 39:27]
  wire  _T_714; // @[LZD.scala 39:25]
  wire [1:0] _T_715; // @[Cat.scala 29:58]
  wire [1:0] _T_716; // @[LZD.scala 44:32]
  wire  _T_717; // @[LZD.scala 39:14]
  wire  _T_718; // @[LZD.scala 39:21]
  wire  _T_719; // @[LZD.scala 39:30]
  wire  _T_720; // @[LZD.scala 39:27]
  wire  _T_721; // @[LZD.scala 39:25]
  wire [1:0] _T_722; // @[Cat.scala 29:58]
  wire  _T_723; // @[Shift.scala 12:21]
  wire  _T_724; // @[Shift.scala 12:21]
  wire  _T_725; // @[LZD.scala 49:16]
  wire  _T_726; // @[LZD.scala 49:27]
  wire  _T_727; // @[LZD.scala 49:25]
  wire  _T_728; // @[LZD.scala 49:47]
  wire  _T_729; // @[LZD.scala 49:59]
  wire  _T_730; // @[LZD.scala 49:35]
  wire [2:0] _T_732; // @[Cat.scala 29:58]
  wire [3:0] _T_733; // @[LZD.scala 44:32]
  wire [1:0] _T_734; // @[LZD.scala 43:32]
  wire  _T_735; // @[LZD.scala 39:14]
  wire  _T_736; // @[LZD.scala 39:21]
  wire  _T_737; // @[LZD.scala 39:30]
  wire  _T_738; // @[LZD.scala 39:27]
  wire  _T_739; // @[LZD.scala 39:25]
  wire [1:0] _T_740; // @[Cat.scala 29:58]
  wire [1:0] _T_741; // @[LZD.scala 44:32]
  wire  _T_742; // @[LZD.scala 39:14]
  wire  _T_743; // @[LZD.scala 39:21]
  wire  _T_744; // @[LZD.scala 39:30]
  wire  _T_745; // @[LZD.scala 39:27]
  wire  _T_746; // @[LZD.scala 39:25]
  wire [1:0] _T_747; // @[Cat.scala 29:58]
  wire  _T_748; // @[Shift.scala 12:21]
  wire  _T_749; // @[Shift.scala 12:21]
  wire  _T_750; // @[LZD.scala 49:16]
  wire  _T_751; // @[LZD.scala 49:27]
  wire  _T_752; // @[LZD.scala 49:25]
  wire  _T_753; // @[LZD.scala 49:47]
  wire  _T_754; // @[LZD.scala 49:59]
  wire  _T_755; // @[LZD.scala 49:35]
  wire [2:0] _T_757; // @[Cat.scala 29:58]
  wire  _T_758; // @[Shift.scala 12:21]
  wire  _T_759; // @[Shift.scala 12:21]
  wire  _T_760; // @[LZD.scala 49:16]
  wire  _T_761; // @[LZD.scala 49:27]
  wire  _T_762; // @[LZD.scala 49:25]
  wire [1:0] _T_763; // @[LZD.scala 49:47]
  wire [1:0] _T_764; // @[LZD.scala 49:59]
  wire [1:0] _T_765; // @[LZD.scala 49:35]
  wire [3:0] _T_767; // @[Cat.scala 29:58]
  wire [1:0] _T_768; // @[LZD.scala 44:32]
  wire  _T_769; // @[LZD.scala 39:14]
  wire  _T_770; // @[LZD.scala 39:21]
  wire  _T_771; // @[LZD.scala 39:30]
  wire  _T_772; // @[LZD.scala 39:27]
  wire  _T_773; // @[LZD.scala 39:25]
  wire  _T_775; // @[Shift.scala 12:21]
  wire [2:0] _T_777; // @[Cat.scala 29:58]
  wire [2:0] _T_778; // @[LZD.scala 55:32]
  wire [2:0] _T_779; // @[LZD.scala 55:20]
  wire [3:0] _T_780; // @[Cat.scala 29:58]
  wire  _T_781; // @[Shift.scala 12:21]
  wire [3:0] _T_783; // @[LZD.scala 55:32]
  wire [3:0] _T_784; // @[LZD.scala 55:20]
  wire [4:0] _T_785; // @[Cat.scala 29:58]
  wire [4:0] _T_786; // @[convert.scala 21:22]
  wire [24:0] _T_787; // @[convert.scala 22:36]
  wire  _T_788; // @[Shift.scala 16:24]
  wire  _T_790; // @[Shift.scala 12:21]
  wire [8:0] _T_791; // @[Shift.scala 64:52]
  wire [24:0] _T_793; // @[Cat.scala 29:58]
  wire [24:0] _T_794; // @[Shift.scala 64:27]
  wire [3:0] _T_795; // @[Shift.scala 66:70]
  wire  _T_796; // @[Shift.scala 12:21]
  wire [16:0] _T_797; // @[Shift.scala 64:52]
  wire [24:0] _T_799; // @[Cat.scala 29:58]
  wire [24:0] _T_800; // @[Shift.scala 64:27]
  wire [2:0] _T_801; // @[Shift.scala 66:70]
  wire  _T_802; // @[Shift.scala 12:21]
  wire [20:0] _T_803; // @[Shift.scala 64:52]
  wire [24:0] _T_805; // @[Cat.scala 29:58]
  wire [24:0] _T_806; // @[Shift.scala 64:27]
  wire [1:0] _T_807; // @[Shift.scala 66:70]
  wire  _T_808; // @[Shift.scala 12:21]
  wire [22:0] _T_809; // @[Shift.scala 64:52]
  wire [24:0] _T_811; // @[Cat.scala 29:58]
  wire [24:0] _T_812; // @[Shift.scala 64:27]
  wire  _T_813; // @[Shift.scala 66:70]
  wire [23:0] _T_815; // @[Shift.scala 64:52]
  wire [24:0] _T_816; // @[Cat.scala 29:58]
  wire [24:0] _T_817; // @[Shift.scala 64:27]
  wire [24:0] _T_818; // @[Shift.scala 16:10]
  wire [2:0] _T_819; // @[convert.scala 23:34]
  wire [21:0] decC_fraction; // @[convert.scala 24:34]
  wire  _T_821; // @[convert.scala 25:26]
  wire [4:0] _T_823; // @[convert.scala 25:42]
  wire [2:0] _T_826; // @[convert.scala 26:67]
  wire [2:0] _T_827; // @[convert.scala 26:51]
  wire [8:0] _T_828; // @[Cat.scala 29:58]
  wire [26:0] _T_830; // @[convert.scala 29:56]
  wire  _T_831; // @[convert.scala 29:60]
  wire  _T_832; // @[convert.scala 29:41]
  wire  decC_isNaR; // @[convert.scala 29:39]
  wire  _T_835; // @[convert.scala 30:19]
  wire  decC_isZero; // @[convert.scala 30:41]
  wire [8:0] decC_scale; // @[convert.scala 32:24]
  wire  _T_843; // @[PositFMA.scala 58:30]
  wire  outIsNaR; // @[PositFMA.scala 58:44]
  wire  _T_844; // @[PositFMA.scala 59:34]
  wire  _T_845; // @[PositFMA.scala 59:47]
  wire  _T_846; // @[PositFMA.scala 59:45]
  wire [23:0] _T_848; // @[Cat.scala 29:58]
  wire [23:0] sigA; // @[PositFMA.scala 59:76]
  wire  _T_849; // @[PositFMA.scala 60:34]
  wire  _T_850; // @[PositFMA.scala 60:47]
  wire  _T_851; // @[PositFMA.scala 60:45]
  wire [23:0] _T_853; // @[Cat.scala 29:58]
  wire [23:0] sigB; // @[PositFMA.scala 60:76]
  wire [47:0] _T_854; // @[PositFMA.scala 61:25]
  wire [47:0] sigP; // @[PositFMA.scala 61:33]
  wire [1:0] head2; // @[PositFMA.scala 62:28]
  wire  _T_855; // @[PositFMA.scala 63:31]
  wire  _T_856; // @[PositFMA.scala 63:25]
  wire  _T_857; // @[PositFMA.scala 63:42]
  wire  addTwo; // @[PositFMA.scala 63:35]
  wire  _T_858; // @[PositFMA.scala 65:23]
  wire  _T_859; // @[PositFMA.scala 65:49]
  wire  addOne; // @[PositFMA.scala 65:43]
  wire [1:0] _T_860; // @[Cat.scala 29:58]
  wire [2:0] expBias; // @[PositFMA.scala 66:39]
  wire  mulSign; // @[PositFMA.scala 67:28]
  wire [9:0] _T_861; // @[PositFMA.scala 69:30]
  wire [9:0] _GEN_12; // @[PositFMA.scala 69:44]
  wire [9:0] _T_863; // @[PositFMA.scala 69:44]
  wire [9:0] mulScale; // @[PositFMA.scala 69:44]
  wire [45:0] _T_864; // @[PositFMA.scala 72:29]
  wire [44:0] _T_865; // @[PositFMA.scala 73:29]
  wire [45:0] _T_866; // @[PositFMA.scala 73:48]
  wire [45:0] mulSigTmp; // @[PositFMA.scala 70:22]
  wire  _T_868; // @[PositFMA.scala 77:39]
  wire  _T_869; // @[PositFMA.scala 77:43]
  wire [44:0] _T_870; // @[PositFMA.scala 78:39]
  wire [46:0] mulSig; // @[Cat.scala 29:58]
  reg  outIsNaR_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg [46:0] mulSig_phase2; // @[Reg.scala 15:16]
  reg [63:0] _RAND_1;
  reg [21:0] addFrac_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [9:0] mulScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [8:0] addScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  addSign_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  addZero_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  inValid_phase2; // @[Valid.scala 117:22]
  reg [31:0] _RAND_7;
  wire  _T_896; // @[PositFMA.scala 107:29]
  wire  _T_897; // @[PositFMA.scala 107:47]
  wire  _T_898; // @[PositFMA.scala 107:45]
  wire [46:0] extAddSig; // @[Cat.scala 29:58]
  wire [9:0] _GEN_13; // @[PositFMA.scala 111:39]
  wire  mulGreater; // @[PositFMA.scala 111:39]
  wire [9:0] greaterScale; // @[PositFMA.scala 112:26]
  wire [9:0] smallerScale; // @[PositFMA.scala 113:26]
  wire [9:0] _T_902; // @[PositFMA.scala 114:36]
  wire [9:0] scaleDiff; // @[PositFMA.scala 114:36]
  wire [46:0] greaterSig; // @[PositFMA.scala 115:26]
  wire [46:0] smallerSigTmp; // @[PositFMA.scala 116:26]
  wire [9:0] _T_903; // @[PositFMA.scala 117:69]
  wire  _T_904; // @[Shift.scala 39:24]
  wire [5:0] _T_905; // @[Shift.scala 40:44]
  wire [14:0] _T_906; // @[Shift.scala 90:30]
  wire [31:0] _T_907; // @[Shift.scala 90:48]
  wire  _T_908; // @[Shift.scala 90:57]
  wire [14:0] _GEN_14; // @[Shift.scala 90:39]
  wire [14:0] _T_909; // @[Shift.scala 90:39]
  wire  _T_910; // @[Shift.scala 12:21]
  wire  _T_911; // @[Shift.scala 12:21]
  wire [31:0] _T_913; // @[Bitwise.scala 71:12]
  wire [46:0] _T_914; // @[Cat.scala 29:58]
  wire [46:0] _T_915; // @[Shift.scala 91:22]
  wire [4:0] _T_916; // @[Shift.scala 92:77]
  wire [30:0] _T_917; // @[Shift.scala 90:30]
  wire [15:0] _T_918; // @[Shift.scala 90:48]
  wire  _T_919; // @[Shift.scala 90:57]
  wire [30:0] _GEN_15; // @[Shift.scala 90:39]
  wire [30:0] _T_920; // @[Shift.scala 90:39]
  wire  _T_921; // @[Shift.scala 12:21]
  wire  _T_922; // @[Shift.scala 12:21]
  wire [15:0] _T_924; // @[Bitwise.scala 71:12]
  wire [46:0] _T_925; // @[Cat.scala 29:58]
  wire [46:0] _T_926; // @[Shift.scala 91:22]
  wire [3:0] _T_927; // @[Shift.scala 92:77]
  wire [38:0] _T_928; // @[Shift.scala 90:30]
  wire [7:0] _T_929; // @[Shift.scala 90:48]
  wire  _T_930; // @[Shift.scala 90:57]
  wire [38:0] _GEN_16; // @[Shift.scala 90:39]
  wire [38:0] _T_931; // @[Shift.scala 90:39]
  wire  _T_932; // @[Shift.scala 12:21]
  wire  _T_933; // @[Shift.scala 12:21]
  wire [7:0] _T_935; // @[Bitwise.scala 71:12]
  wire [46:0] _T_936; // @[Cat.scala 29:58]
  wire [46:0] _T_937; // @[Shift.scala 91:22]
  wire [2:0] _T_938; // @[Shift.scala 92:77]
  wire [42:0] _T_939; // @[Shift.scala 90:30]
  wire [3:0] _T_940; // @[Shift.scala 90:48]
  wire  _T_941; // @[Shift.scala 90:57]
  wire [42:0] _GEN_17; // @[Shift.scala 90:39]
  wire [42:0] _T_942; // @[Shift.scala 90:39]
  wire  _T_943; // @[Shift.scala 12:21]
  wire  _T_944; // @[Shift.scala 12:21]
  wire [3:0] _T_946; // @[Bitwise.scala 71:12]
  wire [46:0] _T_947; // @[Cat.scala 29:58]
  wire [46:0] _T_948; // @[Shift.scala 91:22]
  wire [1:0] _T_949; // @[Shift.scala 92:77]
  wire [44:0] _T_950; // @[Shift.scala 90:30]
  wire [1:0] _T_951; // @[Shift.scala 90:48]
  wire  _T_952; // @[Shift.scala 90:57]
  wire [44:0] _GEN_18; // @[Shift.scala 90:39]
  wire [44:0] _T_953; // @[Shift.scala 90:39]
  wire  _T_954; // @[Shift.scala 12:21]
  wire  _T_955; // @[Shift.scala 12:21]
  wire [1:0] _T_957; // @[Bitwise.scala 71:12]
  wire [46:0] _T_958; // @[Cat.scala 29:58]
  wire [46:0] _T_959; // @[Shift.scala 91:22]
  wire  _T_960; // @[Shift.scala 92:77]
  wire [45:0] _T_961; // @[Shift.scala 90:30]
  wire  _T_962; // @[Shift.scala 90:48]
  wire [45:0] _GEN_19; // @[Shift.scala 90:39]
  wire [45:0] _T_964; // @[Shift.scala 90:39]
  wire  _T_966; // @[Shift.scala 12:21]
  wire [46:0] _T_967; // @[Cat.scala 29:58]
  wire [46:0] _T_968; // @[Shift.scala 91:22]
  wire [46:0] _T_971; // @[Bitwise.scala 71:12]
  wire [46:0] smallerSig; // @[Shift.scala 39:10]
  wire [47:0] rawSumSig; // @[PositFMA.scala 118:34]
  wire  _T_972; // @[PositFMA.scala 119:42]
  wire  _T_973; // @[PositFMA.scala 119:46]
  wire  _T_974; // @[PositFMA.scala 119:79]
  wire  sumSign; // @[PositFMA.scala 119:63]
  wire [46:0] _T_976; // @[PositFMA.scala 120:50]
  wire [47:0] signSumSig; // @[Cat.scala 29:58]
  wire [46:0] _T_977; // @[PositFMA.scala 124:33]
  wire [46:0] _T_978; // @[PositFMA.scala 124:68]
  wire [46:0] sumXor; // @[PositFMA.scala 124:51]
  wire [31:0] _T_979; // @[LZD.scala 43:32]
  wire [15:0] _T_980; // @[LZD.scala 43:32]
  wire [7:0] _T_981; // @[LZD.scala 43:32]
  wire [3:0] _T_982; // @[LZD.scala 43:32]
  wire [1:0] _T_983; // @[LZD.scala 43:32]
  wire  _T_984; // @[LZD.scala 39:14]
  wire  _T_985; // @[LZD.scala 39:21]
  wire  _T_986; // @[LZD.scala 39:30]
  wire  _T_987; // @[LZD.scala 39:27]
  wire  _T_988; // @[LZD.scala 39:25]
  wire [1:0] _T_989; // @[Cat.scala 29:58]
  wire [1:0] _T_990; // @[LZD.scala 44:32]
  wire  _T_991; // @[LZD.scala 39:14]
  wire  _T_992; // @[LZD.scala 39:21]
  wire  _T_993; // @[LZD.scala 39:30]
  wire  _T_994; // @[LZD.scala 39:27]
  wire  _T_995; // @[LZD.scala 39:25]
  wire [1:0] _T_996; // @[Cat.scala 29:58]
  wire  _T_997; // @[Shift.scala 12:21]
  wire  _T_998; // @[Shift.scala 12:21]
  wire  _T_999; // @[LZD.scala 49:16]
  wire  _T_1000; // @[LZD.scala 49:27]
  wire  _T_1001; // @[LZD.scala 49:25]
  wire  _T_1002; // @[LZD.scala 49:47]
  wire  _T_1003; // @[LZD.scala 49:59]
  wire  _T_1004; // @[LZD.scala 49:35]
  wire [2:0] _T_1006; // @[Cat.scala 29:58]
  wire [3:0] _T_1007; // @[LZD.scala 44:32]
  wire [1:0] _T_1008; // @[LZD.scala 43:32]
  wire  _T_1009; // @[LZD.scala 39:14]
  wire  _T_1010; // @[LZD.scala 39:21]
  wire  _T_1011; // @[LZD.scala 39:30]
  wire  _T_1012; // @[LZD.scala 39:27]
  wire  _T_1013; // @[LZD.scala 39:25]
  wire [1:0] _T_1014; // @[Cat.scala 29:58]
  wire [1:0] _T_1015; // @[LZD.scala 44:32]
  wire  _T_1016; // @[LZD.scala 39:14]
  wire  _T_1017; // @[LZD.scala 39:21]
  wire  _T_1018; // @[LZD.scala 39:30]
  wire  _T_1019; // @[LZD.scala 39:27]
  wire  _T_1020; // @[LZD.scala 39:25]
  wire [1:0] _T_1021; // @[Cat.scala 29:58]
  wire  _T_1022; // @[Shift.scala 12:21]
  wire  _T_1023; // @[Shift.scala 12:21]
  wire  _T_1024; // @[LZD.scala 49:16]
  wire  _T_1025; // @[LZD.scala 49:27]
  wire  _T_1026; // @[LZD.scala 49:25]
  wire  _T_1027; // @[LZD.scala 49:47]
  wire  _T_1028; // @[LZD.scala 49:59]
  wire  _T_1029; // @[LZD.scala 49:35]
  wire [2:0] _T_1031; // @[Cat.scala 29:58]
  wire  _T_1032; // @[Shift.scala 12:21]
  wire  _T_1033; // @[Shift.scala 12:21]
  wire  _T_1034; // @[LZD.scala 49:16]
  wire  _T_1035; // @[LZD.scala 49:27]
  wire  _T_1036; // @[LZD.scala 49:25]
  wire [1:0] _T_1037; // @[LZD.scala 49:47]
  wire [1:0] _T_1038; // @[LZD.scala 49:59]
  wire [1:0] _T_1039; // @[LZD.scala 49:35]
  wire [3:0] _T_1041; // @[Cat.scala 29:58]
  wire [7:0] _T_1042; // @[LZD.scala 44:32]
  wire [3:0] _T_1043; // @[LZD.scala 43:32]
  wire [1:0] _T_1044; // @[LZD.scala 43:32]
  wire  _T_1045; // @[LZD.scala 39:14]
  wire  _T_1046; // @[LZD.scala 39:21]
  wire  _T_1047; // @[LZD.scala 39:30]
  wire  _T_1048; // @[LZD.scala 39:27]
  wire  _T_1049; // @[LZD.scala 39:25]
  wire [1:0] _T_1050; // @[Cat.scala 29:58]
  wire [1:0] _T_1051; // @[LZD.scala 44:32]
  wire  _T_1052; // @[LZD.scala 39:14]
  wire  _T_1053; // @[LZD.scala 39:21]
  wire  _T_1054; // @[LZD.scala 39:30]
  wire  _T_1055; // @[LZD.scala 39:27]
  wire  _T_1056; // @[LZD.scala 39:25]
  wire [1:0] _T_1057; // @[Cat.scala 29:58]
  wire  _T_1058; // @[Shift.scala 12:21]
  wire  _T_1059; // @[Shift.scala 12:21]
  wire  _T_1060; // @[LZD.scala 49:16]
  wire  _T_1061; // @[LZD.scala 49:27]
  wire  _T_1062; // @[LZD.scala 49:25]
  wire  _T_1063; // @[LZD.scala 49:47]
  wire  _T_1064; // @[LZD.scala 49:59]
  wire  _T_1065; // @[LZD.scala 49:35]
  wire [2:0] _T_1067; // @[Cat.scala 29:58]
  wire [3:0] _T_1068; // @[LZD.scala 44:32]
  wire [1:0] _T_1069; // @[LZD.scala 43:32]
  wire  _T_1070; // @[LZD.scala 39:14]
  wire  _T_1071; // @[LZD.scala 39:21]
  wire  _T_1072; // @[LZD.scala 39:30]
  wire  _T_1073; // @[LZD.scala 39:27]
  wire  _T_1074; // @[LZD.scala 39:25]
  wire [1:0] _T_1075; // @[Cat.scala 29:58]
  wire [1:0] _T_1076; // @[LZD.scala 44:32]
  wire  _T_1077; // @[LZD.scala 39:14]
  wire  _T_1078; // @[LZD.scala 39:21]
  wire  _T_1079; // @[LZD.scala 39:30]
  wire  _T_1080; // @[LZD.scala 39:27]
  wire  _T_1081; // @[LZD.scala 39:25]
  wire [1:0] _T_1082; // @[Cat.scala 29:58]
  wire  _T_1083; // @[Shift.scala 12:21]
  wire  _T_1084; // @[Shift.scala 12:21]
  wire  _T_1085; // @[LZD.scala 49:16]
  wire  _T_1086; // @[LZD.scala 49:27]
  wire  _T_1087; // @[LZD.scala 49:25]
  wire  _T_1088; // @[LZD.scala 49:47]
  wire  _T_1089; // @[LZD.scala 49:59]
  wire  _T_1090; // @[LZD.scala 49:35]
  wire [2:0] _T_1092; // @[Cat.scala 29:58]
  wire  _T_1093; // @[Shift.scala 12:21]
  wire  _T_1094; // @[Shift.scala 12:21]
  wire  _T_1095; // @[LZD.scala 49:16]
  wire  _T_1096; // @[LZD.scala 49:27]
  wire  _T_1097; // @[LZD.scala 49:25]
  wire [1:0] _T_1098; // @[LZD.scala 49:47]
  wire [1:0] _T_1099; // @[LZD.scala 49:59]
  wire [1:0] _T_1100; // @[LZD.scala 49:35]
  wire [3:0] _T_1102; // @[Cat.scala 29:58]
  wire  _T_1103; // @[Shift.scala 12:21]
  wire  _T_1104; // @[Shift.scala 12:21]
  wire  _T_1105; // @[LZD.scala 49:16]
  wire  _T_1106; // @[LZD.scala 49:27]
  wire  _T_1107; // @[LZD.scala 49:25]
  wire [2:0] _T_1108; // @[LZD.scala 49:47]
  wire [2:0] _T_1109; // @[LZD.scala 49:59]
  wire [2:0] _T_1110; // @[LZD.scala 49:35]
  wire [4:0] _T_1112; // @[Cat.scala 29:58]
  wire [15:0] _T_1113; // @[LZD.scala 44:32]
  wire [7:0] _T_1114; // @[LZD.scala 43:32]
  wire [3:0] _T_1115; // @[LZD.scala 43:32]
  wire [1:0] _T_1116; // @[LZD.scala 43:32]
  wire  _T_1117; // @[LZD.scala 39:14]
  wire  _T_1118; // @[LZD.scala 39:21]
  wire  _T_1119; // @[LZD.scala 39:30]
  wire  _T_1120; // @[LZD.scala 39:27]
  wire  _T_1121; // @[LZD.scala 39:25]
  wire [1:0] _T_1122; // @[Cat.scala 29:58]
  wire [1:0] _T_1123; // @[LZD.scala 44:32]
  wire  _T_1124; // @[LZD.scala 39:14]
  wire  _T_1125; // @[LZD.scala 39:21]
  wire  _T_1126; // @[LZD.scala 39:30]
  wire  _T_1127; // @[LZD.scala 39:27]
  wire  _T_1128; // @[LZD.scala 39:25]
  wire [1:0] _T_1129; // @[Cat.scala 29:58]
  wire  _T_1130; // @[Shift.scala 12:21]
  wire  _T_1131; // @[Shift.scala 12:21]
  wire  _T_1132; // @[LZD.scala 49:16]
  wire  _T_1133; // @[LZD.scala 49:27]
  wire  _T_1134; // @[LZD.scala 49:25]
  wire  _T_1135; // @[LZD.scala 49:47]
  wire  _T_1136; // @[LZD.scala 49:59]
  wire  _T_1137; // @[LZD.scala 49:35]
  wire [2:0] _T_1139; // @[Cat.scala 29:58]
  wire [3:0] _T_1140; // @[LZD.scala 44:32]
  wire [1:0] _T_1141; // @[LZD.scala 43:32]
  wire  _T_1142; // @[LZD.scala 39:14]
  wire  _T_1143; // @[LZD.scala 39:21]
  wire  _T_1144; // @[LZD.scala 39:30]
  wire  _T_1145; // @[LZD.scala 39:27]
  wire  _T_1146; // @[LZD.scala 39:25]
  wire [1:0] _T_1147; // @[Cat.scala 29:58]
  wire [1:0] _T_1148; // @[LZD.scala 44:32]
  wire  _T_1149; // @[LZD.scala 39:14]
  wire  _T_1150; // @[LZD.scala 39:21]
  wire  _T_1151; // @[LZD.scala 39:30]
  wire  _T_1152; // @[LZD.scala 39:27]
  wire  _T_1153; // @[LZD.scala 39:25]
  wire [1:0] _T_1154; // @[Cat.scala 29:58]
  wire  _T_1155; // @[Shift.scala 12:21]
  wire  _T_1156; // @[Shift.scala 12:21]
  wire  _T_1157; // @[LZD.scala 49:16]
  wire  _T_1158; // @[LZD.scala 49:27]
  wire  _T_1159; // @[LZD.scala 49:25]
  wire  _T_1160; // @[LZD.scala 49:47]
  wire  _T_1161; // @[LZD.scala 49:59]
  wire  _T_1162; // @[LZD.scala 49:35]
  wire [2:0] _T_1164; // @[Cat.scala 29:58]
  wire  _T_1165; // @[Shift.scala 12:21]
  wire  _T_1166; // @[Shift.scala 12:21]
  wire  _T_1167; // @[LZD.scala 49:16]
  wire  _T_1168; // @[LZD.scala 49:27]
  wire  _T_1169; // @[LZD.scala 49:25]
  wire [1:0] _T_1170; // @[LZD.scala 49:47]
  wire [1:0] _T_1171; // @[LZD.scala 49:59]
  wire [1:0] _T_1172; // @[LZD.scala 49:35]
  wire [3:0] _T_1174; // @[Cat.scala 29:58]
  wire [7:0] _T_1175; // @[LZD.scala 44:32]
  wire [3:0] _T_1176; // @[LZD.scala 43:32]
  wire [1:0] _T_1177; // @[LZD.scala 43:32]
  wire  _T_1178; // @[LZD.scala 39:14]
  wire  _T_1179; // @[LZD.scala 39:21]
  wire  _T_1180; // @[LZD.scala 39:30]
  wire  _T_1181; // @[LZD.scala 39:27]
  wire  _T_1182; // @[LZD.scala 39:25]
  wire [1:0] _T_1183; // @[Cat.scala 29:58]
  wire [1:0] _T_1184; // @[LZD.scala 44:32]
  wire  _T_1185; // @[LZD.scala 39:14]
  wire  _T_1186; // @[LZD.scala 39:21]
  wire  _T_1187; // @[LZD.scala 39:30]
  wire  _T_1188; // @[LZD.scala 39:27]
  wire  _T_1189; // @[LZD.scala 39:25]
  wire [1:0] _T_1190; // @[Cat.scala 29:58]
  wire  _T_1191; // @[Shift.scala 12:21]
  wire  _T_1192; // @[Shift.scala 12:21]
  wire  _T_1193; // @[LZD.scala 49:16]
  wire  _T_1194; // @[LZD.scala 49:27]
  wire  _T_1195; // @[LZD.scala 49:25]
  wire  _T_1196; // @[LZD.scala 49:47]
  wire  _T_1197; // @[LZD.scala 49:59]
  wire  _T_1198; // @[LZD.scala 49:35]
  wire [2:0] _T_1200; // @[Cat.scala 29:58]
  wire [3:0] _T_1201; // @[LZD.scala 44:32]
  wire [1:0] _T_1202; // @[LZD.scala 43:32]
  wire  _T_1203; // @[LZD.scala 39:14]
  wire  _T_1204; // @[LZD.scala 39:21]
  wire  _T_1205; // @[LZD.scala 39:30]
  wire  _T_1206; // @[LZD.scala 39:27]
  wire  _T_1207; // @[LZD.scala 39:25]
  wire [1:0] _T_1208; // @[Cat.scala 29:58]
  wire [1:0] _T_1209; // @[LZD.scala 44:32]
  wire  _T_1210; // @[LZD.scala 39:14]
  wire  _T_1211; // @[LZD.scala 39:21]
  wire  _T_1212; // @[LZD.scala 39:30]
  wire  _T_1213; // @[LZD.scala 39:27]
  wire  _T_1214; // @[LZD.scala 39:25]
  wire [1:0] _T_1215; // @[Cat.scala 29:58]
  wire  _T_1216; // @[Shift.scala 12:21]
  wire  _T_1217; // @[Shift.scala 12:21]
  wire  _T_1218; // @[LZD.scala 49:16]
  wire  _T_1219; // @[LZD.scala 49:27]
  wire  _T_1220; // @[LZD.scala 49:25]
  wire  _T_1221; // @[LZD.scala 49:47]
  wire  _T_1222; // @[LZD.scala 49:59]
  wire  _T_1223; // @[LZD.scala 49:35]
  wire [2:0] _T_1225; // @[Cat.scala 29:58]
  wire  _T_1226; // @[Shift.scala 12:21]
  wire  _T_1227; // @[Shift.scala 12:21]
  wire  _T_1228; // @[LZD.scala 49:16]
  wire  _T_1229; // @[LZD.scala 49:27]
  wire  _T_1230; // @[LZD.scala 49:25]
  wire [1:0] _T_1231; // @[LZD.scala 49:47]
  wire [1:0] _T_1232; // @[LZD.scala 49:59]
  wire [1:0] _T_1233; // @[LZD.scala 49:35]
  wire [3:0] _T_1235; // @[Cat.scala 29:58]
  wire  _T_1236; // @[Shift.scala 12:21]
  wire  _T_1237; // @[Shift.scala 12:21]
  wire  _T_1238; // @[LZD.scala 49:16]
  wire  _T_1239; // @[LZD.scala 49:27]
  wire  _T_1240; // @[LZD.scala 49:25]
  wire [2:0] _T_1241; // @[LZD.scala 49:47]
  wire [2:0] _T_1242; // @[LZD.scala 49:59]
  wire [2:0] _T_1243; // @[LZD.scala 49:35]
  wire [4:0] _T_1245; // @[Cat.scala 29:58]
  wire  _T_1246; // @[Shift.scala 12:21]
  wire  _T_1247; // @[Shift.scala 12:21]
  wire  _T_1248; // @[LZD.scala 49:16]
  wire  _T_1249; // @[LZD.scala 49:27]
  wire  _T_1250; // @[LZD.scala 49:25]
  wire [3:0] _T_1251; // @[LZD.scala 49:47]
  wire [3:0] _T_1252; // @[LZD.scala 49:59]
  wire [3:0] _T_1253; // @[LZD.scala 49:35]
  wire [5:0] _T_1255; // @[Cat.scala 29:58]
  wire [14:0] _T_1256; // @[LZD.scala 44:32]
  wire [7:0] _T_1257; // @[LZD.scala 43:32]
  wire [3:0] _T_1258; // @[LZD.scala 43:32]
  wire [1:0] _T_1259; // @[LZD.scala 43:32]
  wire  _T_1260; // @[LZD.scala 39:14]
  wire  _T_1261; // @[LZD.scala 39:21]
  wire  _T_1262; // @[LZD.scala 39:30]
  wire  _T_1263; // @[LZD.scala 39:27]
  wire  _T_1264; // @[LZD.scala 39:25]
  wire [1:0] _T_1265; // @[Cat.scala 29:58]
  wire [1:0] _T_1266; // @[LZD.scala 44:32]
  wire  _T_1267; // @[LZD.scala 39:14]
  wire  _T_1268; // @[LZD.scala 39:21]
  wire  _T_1269; // @[LZD.scala 39:30]
  wire  _T_1270; // @[LZD.scala 39:27]
  wire  _T_1271; // @[LZD.scala 39:25]
  wire [1:0] _T_1272; // @[Cat.scala 29:58]
  wire  _T_1273; // @[Shift.scala 12:21]
  wire  _T_1274; // @[Shift.scala 12:21]
  wire  _T_1275; // @[LZD.scala 49:16]
  wire  _T_1276; // @[LZD.scala 49:27]
  wire  _T_1277; // @[LZD.scala 49:25]
  wire  _T_1278; // @[LZD.scala 49:47]
  wire  _T_1279; // @[LZD.scala 49:59]
  wire  _T_1280; // @[LZD.scala 49:35]
  wire [2:0] _T_1282; // @[Cat.scala 29:58]
  wire [3:0] _T_1283; // @[LZD.scala 44:32]
  wire [1:0] _T_1284; // @[LZD.scala 43:32]
  wire  _T_1285; // @[LZD.scala 39:14]
  wire  _T_1286; // @[LZD.scala 39:21]
  wire  _T_1287; // @[LZD.scala 39:30]
  wire  _T_1288; // @[LZD.scala 39:27]
  wire  _T_1289; // @[LZD.scala 39:25]
  wire [1:0] _T_1290; // @[Cat.scala 29:58]
  wire [1:0] _T_1291; // @[LZD.scala 44:32]
  wire  _T_1292; // @[LZD.scala 39:14]
  wire  _T_1293; // @[LZD.scala 39:21]
  wire  _T_1294; // @[LZD.scala 39:30]
  wire  _T_1295; // @[LZD.scala 39:27]
  wire  _T_1296; // @[LZD.scala 39:25]
  wire [1:0] _T_1297; // @[Cat.scala 29:58]
  wire  _T_1298; // @[Shift.scala 12:21]
  wire  _T_1299; // @[Shift.scala 12:21]
  wire  _T_1300; // @[LZD.scala 49:16]
  wire  _T_1301; // @[LZD.scala 49:27]
  wire  _T_1302; // @[LZD.scala 49:25]
  wire  _T_1303; // @[LZD.scala 49:47]
  wire  _T_1304; // @[LZD.scala 49:59]
  wire  _T_1305; // @[LZD.scala 49:35]
  wire [2:0] _T_1307; // @[Cat.scala 29:58]
  wire  _T_1308; // @[Shift.scala 12:21]
  wire  _T_1309; // @[Shift.scala 12:21]
  wire  _T_1310; // @[LZD.scala 49:16]
  wire  _T_1311; // @[LZD.scala 49:27]
  wire  _T_1312; // @[LZD.scala 49:25]
  wire [1:0] _T_1313; // @[LZD.scala 49:47]
  wire [1:0] _T_1314; // @[LZD.scala 49:59]
  wire [1:0] _T_1315; // @[LZD.scala 49:35]
  wire [3:0] _T_1317; // @[Cat.scala 29:58]
  wire [6:0] _T_1318; // @[LZD.scala 44:32]
  wire [3:0] _T_1319; // @[LZD.scala 43:32]
  wire [1:0] _T_1320; // @[LZD.scala 43:32]
  wire  _T_1321; // @[LZD.scala 39:14]
  wire  _T_1322; // @[LZD.scala 39:21]
  wire  _T_1323; // @[LZD.scala 39:30]
  wire  _T_1324; // @[LZD.scala 39:27]
  wire  _T_1325; // @[LZD.scala 39:25]
  wire [1:0] _T_1326; // @[Cat.scala 29:58]
  wire [1:0] _T_1327; // @[LZD.scala 44:32]
  wire  _T_1328; // @[LZD.scala 39:14]
  wire  _T_1329; // @[LZD.scala 39:21]
  wire  _T_1330; // @[LZD.scala 39:30]
  wire  _T_1331; // @[LZD.scala 39:27]
  wire  _T_1332; // @[LZD.scala 39:25]
  wire [1:0] _T_1333; // @[Cat.scala 29:58]
  wire  _T_1334; // @[Shift.scala 12:21]
  wire  _T_1335; // @[Shift.scala 12:21]
  wire  _T_1336; // @[LZD.scala 49:16]
  wire  _T_1337; // @[LZD.scala 49:27]
  wire  _T_1338; // @[LZD.scala 49:25]
  wire  _T_1339; // @[LZD.scala 49:47]
  wire  _T_1340; // @[LZD.scala 49:59]
  wire  _T_1341; // @[LZD.scala 49:35]
  wire [2:0] _T_1343; // @[Cat.scala 29:58]
  wire [2:0] _T_1344; // @[LZD.scala 44:32]
  wire [1:0] _T_1345; // @[LZD.scala 43:32]
  wire  _T_1346; // @[LZD.scala 39:14]
  wire  _T_1347; // @[LZD.scala 39:21]
  wire  _T_1348; // @[LZD.scala 39:30]
  wire  _T_1349; // @[LZD.scala 39:27]
  wire  _T_1350; // @[LZD.scala 39:25]
  wire [1:0] _T_1351; // @[Cat.scala 29:58]
  wire  _T_1352; // @[LZD.scala 44:32]
  wire  _T_1354; // @[Shift.scala 12:21]
  wire  _T_1356; // @[LZD.scala 55:32]
  wire  _T_1357; // @[LZD.scala 55:20]
  wire [1:0] _T_1358; // @[Cat.scala 29:58]
  wire  _T_1359; // @[Shift.scala 12:21]
  wire [1:0] _T_1361; // @[LZD.scala 55:32]
  wire [1:0] _T_1362; // @[LZD.scala 55:20]
  wire [2:0] _T_1363; // @[Cat.scala 29:58]
  wire  _T_1364; // @[Shift.scala 12:21]
  wire [2:0] _T_1366; // @[LZD.scala 55:32]
  wire [2:0] _T_1367; // @[LZD.scala 55:20]
  wire  _T_1369; // @[Shift.scala 12:21]
  wire [4:0] _T_1371; // @[Cat.scala 29:58]
  wire [4:0] _T_1372; // @[LZD.scala 55:32]
  wire [4:0] _T_1373; // @[LZD.scala 55:20]
  wire [5:0] sumLZD; // @[Cat.scala 29:58]
  wire [5:0] shiftValue; // @[PositFMA.scala 126:24]
  wire [45:0] _T_1374; // @[PositFMA.scala 127:38]
  wire  _T_1375; // @[Shift.scala 16:24]
  wire  _T_1377; // @[Shift.scala 12:21]
  wire [13:0] _T_1378; // @[Shift.scala 64:52]
  wire [45:0] _T_1380; // @[Cat.scala 29:58]
  wire [45:0] _T_1381; // @[Shift.scala 64:27]
  wire [4:0] _T_1382; // @[Shift.scala 66:70]
  wire  _T_1383; // @[Shift.scala 12:21]
  wire [29:0] _T_1384; // @[Shift.scala 64:52]
  wire [45:0] _T_1386; // @[Cat.scala 29:58]
  wire [45:0] _T_1387; // @[Shift.scala 64:27]
  wire [3:0] _T_1388; // @[Shift.scala 66:70]
  wire  _T_1389; // @[Shift.scala 12:21]
  wire [37:0] _T_1390; // @[Shift.scala 64:52]
  wire [45:0] _T_1392; // @[Cat.scala 29:58]
  wire [45:0] _T_1393; // @[Shift.scala 64:27]
  wire [2:0] _T_1394; // @[Shift.scala 66:70]
  wire  _T_1395; // @[Shift.scala 12:21]
  wire [41:0] _T_1396; // @[Shift.scala 64:52]
  wire [45:0] _T_1398; // @[Cat.scala 29:58]
  wire [45:0] _T_1399; // @[Shift.scala 64:27]
  wire [1:0] _T_1400; // @[Shift.scala 66:70]
  wire  _T_1401; // @[Shift.scala 12:21]
  wire [43:0] _T_1402; // @[Shift.scala 64:52]
  wire [45:0] _T_1404; // @[Cat.scala 29:58]
  wire [45:0] _T_1405; // @[Shift.scala 64:27]
  wire  _T_1406; // @[Shift.scala 66:70]
  wire [44:0] _T_1408; // @[Shift.scala 64:52]
  wire [45:0] _T_1409; // @[Cat.scala 29:58]
  wire [45:0] _T_1410; // @[Shift.scala 64:27]
  wire [45:0] normalFracTmp; // @[Shift.scala 16:10]
  wire [9:0] _T_1412; // @[PositFMA.scala 130:36]
  wire [9:0] _T_1413; // @[PositFMA.scala 130:36]
  wire [6:0] _T_1414; // @[Cat.scala 29:58]
  wire [6:0] _T_1415; // @[PositFMA.scala 130:61]
  wire [9:0] _GEN_20; // @[PositFMA.scala 130:42]
  wire [9:0] _T_1417; // @[PositFMA.scala 130:42]
  wire [9:0] sumScale; // @[PositFMA.scala 130:42]
  wire [21:0] sumFrac; // @[PositFMA.scala 131:41]
  wire [23:0] grsTmp; // @[PositFMA.scala 134:41]
  wire [1:0] _T_1418; // @[PositFMA.scala 137:40]
  wire [21:0] _T_1419; // @[PositFMA.scala 137:56]
  wire  _T_1420; // @[PositFMA.scala 137:60]
  wire  underflow; // @[PositFMA.scala 144:32]
  wire  overflow; // @[PositFMA.scala 145:32]
  wire  _T_1421; // @[PositFMA.scala 154:32]
  wire  decF_isZero; // @[PositFMA.scala 154:20]
  wire [9:0] _T_1423; // @[Mux.scala 87:16]
  wire [9:0] _T_1424; // @[Mux.scala 87:16]
  wire [8:0] _GEN_21; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  wire [8:0] decF_scale; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  wire [2:0] _T_1425; // @[convert.scala 46:61]
  wire [2:0] _T_1426; // @[convert.scala 46:52]
  wire [2:0] _T_1428; // @[convert.scala 46:42]
  wire [5:0] _T_1429; // @[convert.scala 48:34]
  wire  _T_1430; // @[convert.scala 49:36]
  wire [5:0] _T_1432; // @[convert.scala 50:36]
  wire [5:0] _T_1433; // @[convert.scala 50:36]
  wire [5:0] _T_1434; // @[convert.scala 50:28]
  wire  _T_1435; // @[convert.scala 51:31]
  wire  _T_1436; // @[convert.scala 52:43]
  wire [29:0] _T_1440; // @[Cat.scala 29:58]
  wire [5:0] _T_1441; // @[Shift.scala 39:17]
  wire  _T_1442; // @[Shift.scala 39:24]
  wire [4:0] _T_1443; // @[Shift.scala 40:44]
  wire [13:0] _T_1444; // @[Shift.scala 90:30]
  wire [15:0] _T_1445; // @[Shift.scala 90:48]
  wire  _T_1446; // @[Shift.scala 90:57]
  wire [13:0] _GEN_22; // @[Shift.scala 90:39]
  wire [13:0] _T_1447; // @[Shift.scala 90:39]
  wire  _T_1448; // @[Shift.scala 12:21]
  wire  _T_1449; // @[Shift.scala 12:21]
  wire [15:0] _T_1451; // @[Bitwise.scala 71:12]
  wire [29:0] _T_1452; // @[Cat.scala 29:58]
  wire [29:0] _T_1453; // @[Shift.scala 91:22]
  wire [3:0] _T_1454; // @[Shift.scala 92:77]
  wire [21:0] _T_1455; // @[Shift.scala 90:30]
  wire [7:0] _T_1456; // @[Shift.scala 90:48]
  wire  _T_1457; // @[Shift.scala 90:57]
  wire [21:0] _GEN_23; // @[Shift.scala 90:39]
  wire [21:0] _T_1458; // @[Shift.scala 90:39]
  wire  _T_1459; // @[Shift.scala 12:21]
  wire  _T_1460; // @[Shift.scala 12:21]
  wire [7:0] _T_1462; // @[Bitwise.scala 71:12]
  wire [29:0] _T_1463; // @[Cat.scala 29:58]
  wire [29:0] _T_1464; // @[Shift.scala 91:22]
  wire [2:0] _T_1465; // @[Shift.scala 92:77]
  wire [25:0] _T_1466; // @[Shift.scala 90:30]
  wire [3:0] _T_1467; // @[Shift.scala 90:48]
  wire  _T_1468; // @[Shift.scala 90:57]
  wire [25:0] _GEN_24; // @[Shift.scala 90:39]
  wire [25:0] _T_1469; // @[Shift.scala 90:39]
  wire  _T_1470; // @[Shift.scala 12:21]
  wire  _T_1471; // @[Shift.scala 12:21]
  wire [3:0] _T_1473; // @[Bitwise.scala 71:12]
  wire [29:0] _T_1474; // @[Cat.scala 29:58]
  wire [29:0] _T_1475; // @[Shift.scala 91:22]
  wire [1:0] _T_1476; // @[Shift.scala 92:77]
  wire [27:0] _T_1477; // @[Shift.scala 90:30]
  wire [1:0] _T_1478; // @[Shift.scala 90:48]
  wire  _T_1479; // @[Shift.scala 90:57]
  wire [27:0] _GEN_25; // @[Shift.scala 90:39]
  wire [27:0] _T_1480; // @[Shift.scala 90:39]
  wire  _T_1481; // @[Shift.scala 12:21]
  wire  _T_1482; // @[Shift.scala 12:21]
  wire [1:0] _T_1484; // @[Bitwise.scala 71:12]
  wire [29:0] _T_1485; // @[Cat.scala 29:58]
  wire [29:0] _T_1486; // @[Shift.scala 91:22]
  wire  _T_1487; // @[Shift.scala 92:77]
  wire [28:0] _T_1488; // @[Shift.scala 90:30]
  wire  _T_1489; // @[Shift.scala 90:48]
  wire [28:0] _GEN_26; // @[Shift.scala 90:39]
  wire [28:0] _T_1491; // @[Shift.scala 90:39]
  wire  _T_1493; // @[Shift.scala 12:21]
  wire [29:0] _T_1494; // @[Cat.scala 29:58]
  wire [29:0] _T_1495; // @[Shift.scala 91:22]
  wire [29:0] _T_1498; // @[Bitwise.scala 71:12]
  wire [29:0] _T_1499; // @[Shift.scala 39:10]
  wire  _T_1500; // @[convert.scala 55:31]
  wire  _T_1501; // @[convert.scala 56:31]
  wire  _T_1502; // @[convert.scala 57:31]
  wire  _T_1503; // @[convert.scala 58:31]
  wire [26:0] _T_1504; // @[convert.scala 59:69]
  wire  _T_1505; // @[convert.scala 59:81]
  wire  _T_1506; // @[convert.scala 59:50]
  wire  _T_1508; // @[convert.scala 60:81]
  wire  _T_1509; // @[convert.scala 61:44]
  wire  _T_1510; // @[convert.scala 61:52]
  wire  _T_1511; // @[convert.scala 61:36]
  wire  _T_1512; // @[convert.scala 62:63]
  wire  _T_1513; // @[convert.scala 62:103]
  wire  _T_1514; // @[convert.scala 62:60]
  wire [26:0] _GEN_27; // @[convert.scala 63:56]
  wire [26:0] _T_1517; // @[convert.scala 63:56]
  wire [27:0] _T_1518; // @[Cat.scala 29:58]
  reg  _T_1522; // @[Valid.scala 117:22]
  reg [31:0] _RAND_8;
  reg [27:0] _T_1526; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  assign _T = io_fmaOp[1]; // @[PositFMA.scala 47:36]
  assign _T_2 = _T ? 28'hfffffff : 28'h0; // @[Bitwise.scala 71:12]
  assign _T_3 = _T_2 ^ io_A; // @[PositFMA.scala 47:41]
  assign _GEN_10 = {{27'd0}, _T}; // @[PositFMA.scala 47:49]
  assign realA = _T_3 + _GEN_10; // @[PositFMA.scala 47:49]
  assign _T_6 = io_fmaOp[0]; // @[PositFMA.scala 48:36]
  assign _T_8 = _T_6 ? 28'hfffffff : 28'h0; // @[Bitwise.scala 71:12]
  assign _T_9 = _T_8 ^ io_C; // @[PositFMA.scala 48:41]
  assign _GEN_11 = {{27'd0}, _T_6}; // @[PositFMA.scala 48:49]
  assign realC = _T_9 + _GEN_11; // @[PositFMA.scala 48:49]
  assign _T_13 = realA[27]; // @[convert.scala 18:24]
  assign _T_14 = realA[26]; // @[convert.scala 18:40]
  assign _T_15 = _T_13 ^ _T_14; // @[convert.scala 18:36]
  assign _T_16 = realA[26:1]; // @[convert.scala 19:24]
  assign _T_17 = realA[25:0]; // @[convert.scala 19:43]
  assign _T_18 = _T_16 ^ _T_17; // @[convert.scala 19:39]
  assign _T_19 = _T_18[25:10]; // @[LZD.scala 43:32]
  assign _T_20 = _T_19[15:8]; // @[LZD.scala 43:32]
  assign _T_21 = _T_20[7:4]; // @[LZD.scala 43:32]
  assign _T_22 = _T_21[3:2]; // @[LZD.scala 43:32]
  assign _T_23 = _T_22 != 2'h0; // @[LZD.scala 39:14]
  assign _T_24 = _T_22[1]; // @[LZD.scala 39:21]
  assign _T_25 = _T_22[0]; // @[LZD.scala 39:30]
  assign _T_26 = ~ _T_25; // @[LZD.scala 39:27]
  assign _T_27 = _T_24 | _T_26; // @[LZD.scala 39:25]
  assign _T_28 = {_T_23,_T_27}; // @[Cat.scala 29:58]
  assign _T_29 = _T_21[1:0]; // @[LZD.scala 44:32]
  assign _T_30 = _T_29 != 2'h0; // @[LZD.scala 39:14]
  assign _T_31 = _T_29[1]; // @[LZD.scala 39:21]
  assign _T_32 = _T_29[0]; // @[LZD.scala 39:30]
  assign _T_33 = ~ _T_32; // @[LZD.scala 39:27]
  assign _T_34 = _T_31 | _T_33; // @[LZD.scala 39:25]
  assign _T_35 = {_T_30,_T_34}; // @[Cat.scala 29:58]
  assign _T_36 = _T_28[1]; // @[Shift.scala 12:21]
  assign _T_37 = _T_35[1]; // @[Shift.scala 12:21]
  assign _T_38 = _T_36 | _T_37; // @[LZD.scala 49:16]
  assign _T_39 = ~ _T_37; // @[LZD.scala 49:27]
  assign _T_40 = _T_36 | _T_39; // @[LZD.scala 49:25]
  assign _T_41 = _T_28[0:0]; // @[LZD.scala 49:47]
  assign _T_42 = _T_35[0:0]; // @[LZD.scala 49:59]
  assign _T_43 = _T_36 ? _T_41 : _T_42; // @[LZD.scala 49:35]
  assign _T_45 = {_T_38,_T_40,_T_43}; // @[Cat.scala 29:58]
  assign _T_46 = _T_20[3:0]; // @[LZD.scala 44:32]
  assign _T_47 = _T_46[3:2]; // @[LZD.scala 43:32]
  assign _T_48 = _T_47 != 2'h0; // @[LZD.scala 39:14]
  assign _T_49 = _T_47[1]; // @[LZD.scala 39:21]
  assign _T_50 = _T_47[0]; // @[LZD.scala 39:30]
  assign _T_51 = ~ _T_50; // @[LZD.scala 39:27]
  assign _T_52 = _T_49 | _T_51; // @[LZD.scala 39:25]
  assign _T_53 = {_T_48,_T_52}; // @[Cat.scala 29:58]
  assign _T_54 = _T_46[1:0]; // @[LZD.scala 44:32]
  assign _T_55 = _T_54 != 2'h0; // @[LZD.scala 39:14]
  assign _T_56 = _T_54[1]; // @[LZD.scala 39:21]
  assign _T_57 = _T_54[0]; // @[LZD.scala 39:30]
  assign _T_58 = ~ _T_57; // @[LZD.scala 39:27]
  assign _T_59 = _T_56 | _T_58; // @[LZD.scala 39:25]
  assign _T_60 = {_T_55,_T_59}; // @[Cat.scala 29:58]
  assign _T_61 = _T_53[1]; // @[Shift.scala 12:21]
  assign _T_62 = _T_60[1]; // @[Shift.scala 12:21]
  assign _T_63 = _T_61 | _T_62; // @[LZD.scala 49:16]
  assign _T_64 = ~ _T_62; // @[LZD.scala 49:27]
  assign _T_65 = _T_61 | _T_64; // @[LZD.scala 49:25]
  assign _T_66 = _T_53[0:0]; // @[LZD.scala 49:47]
  assign _T_67 = _T_60[0:0]; // @[LZD.scala 49:59]
  assign _T_68 = _T_61 ? _T_66 : _T_67; // @[LZD.scala 49:35]
  assign _T_70 = {_T_63,_T_65,_T_68}; // @[Cat.scala 29:58]
  assign _T_71 = _T_45[2]; // @[Shift.scala 12:21]
  assign _T_72 = _T_70[2]; // @[Shift.scala 12:21]
  assign _T_73 = _T_71 | _T_72; // @[LZD.scala 49:16]
  assign _T_74 = ~ _T_72; // @[LZD.scala 49:27]
  assign _T_75 = _T_71 | _T_74; // @[LZD.scala 49:25]
  assign _T_76 = _T_45[1:0]; // @[LZD.scala 49:47]
  assign _T_77 = _T_70[1:0]; // @[LZD.scala 49:59]
  assign _T_78 = _T_71 ? _T_76 : _T_77; // @[LZD.scala 49:35]
  assign _T_80 = {_T_73,_T_75,_T_78}; // @[Cat.scala 29:58]
  assign _T_81 = _T_19[7:0]; // @[LZD.scala 44:32]
  assign _T_82 = _T_81[7:4]; // @[LZD.scala 43:32]
  assign _T_83 = _T_82[3:2]; // @[LZD.scala 43:32]
  assign _T_84 = _T_83 != 2'h0; // @[LZD.scala 39:14]
  assign _T_85 = _T_83[1]; // @[LZD.scala 39:21]
  assign _T_86 = _T_83[0]; // @[LZD.scala 39:30]
  assign _T_87 = ~ _T_86; // @[LZD.scala 39:27]
  assign _T_88 = _T_85 | _T_87; // @[LZD.scala 39:25]
  assign _T_89 = {_T_84,_T_88}; // @[Cat.scala 29:58]
  assign _T_90 = _T_82[1:0]; // @[LZD.scala 44:32]
  assign _T_91 = _T_90 != 2'h0; // @[LZD.scala 39:14]
  assign _T_92 = _T_90[1]; // @[LZD.scala 39:21]
  assign _T_93 = _T_90[0]; // @[LZD.scala 39:30]
  assign _T_94 = ~ _T_93; // @[LZD.scala 39:27]
  assign _T_95 = _T_92 | _T_94; // @[LZD.scala 39:25]
  assign _T_96 = {_T_91,_T_95}; // @[Cat.scala 29:58]
  assign _T_97 = _T_89[1]; // @[Shift.scala 12:21]
  assign _T_98 = _T_96[1]; // @[Shift.scala 12:21]
  assign _T_99 = _T_97 | _T_98; // @[LZD.scala 49:16]
  assign _T_100 = ~ _T_98; // @[LZD.scala 49:27]
  assign _T_101 = _T_97 | _T_100; // @[LZD.scala 49:25]
  assign _T_102 = _T_89[0:0]; // @[LZD.scala 49:47]
  assign _T_103 = _T_96[0:0]; // @[LZD.scala 49:59]
  assign _T_104 = _T_97 ? _T_102 : _T_103; // @[LZD.scala 49:35]
  assign _T_106 = {_T_99,_T_101,_T_104}; // @[Cat.scala 29:58]
  assign _T_107 = _T_81[3:0]; // @[LZD.scala 44:32]
  assign _T_108 = _T_107[3:2]; // @[LZD.scala 43:32]
  assign _T_109 = _T_108 != 2'h0; // @[LZD.scala 39:14]
  assign _T_110 = _T_108[1]; // @[LZD.scala 39:21]
  assign _T_111 = _T_108[0]; // @[LZD.scala 39:30]
  assign _T_112 = ~ _T_111; // @[LZD.scala 39:27]
  assign _T_113 = _T_110 | _T_112; // @[LZD.scala 39:25]
  assign _T_114 = {_T_109,_T_113}; // @[Cat.scala 29:58]
  assign _T_115 = _T_107[1:0]; // @[LZD.scala 44:32]
  assign _T_116 = _T_115 != 2'h0; // @[LZD.scala 39:14]
  assign _T_117 = _T_115[1]; // @[LZD.scala 39:21]
  assign _T_118 = _T_115[0]; // @[LZD.scala 39:30]
  assign _T_119 = ~ _T_118; // @[LZD.scala 39:27]
  assign _T_120 = _T_117 | _T_119; // @[LZD.scala 39:25]
  assign _T_121 = {_T_116,_T_120}; // @[Cat.scala 29:58]
  assign _T_122 = _T_114[1]; // @[Shift.scala 12:21]
  assign _T_123 = _T_121[1]; // @[Shift.scala 12:21]
  assign _T_124 = _T_122 | _T_123; // @[LZD.scala 49:16]
  assign _T_125 = ~ _T_123; // @[LZD.scala 49:27]
  assign _T_126 = _T_122 | _T_125; // @[LZD.scala 49:25]
  assign _T_127 = _T_114[0:0]; // @[LZD.scala 49:47]
  assign _T_128 = _T_121[0:0]; // @[LZD.scala 49:59]
  assign _T_129 = _T_122 ? _T_127 : _T_128; // @[LZD.scala 49:35]
  assign _T_131 = {_T_124,_T_126,_T_129}; // @[Cat.scala 29:58]
  assign _T_132 = _T_106[2]; // @[Shift.scala 12:21]
  assign _T_133 = _T_131[2]; // @[Shift.scala 12:21]
  assign _T_134 = _T_132 | _T_133; // @[LZD.scala 49:16]
  assign _T_135 = ~ _T_133; // @[LZD.scala 49:27]
  assign _T_136 = _T_132 | _T_135; // @[LZD.scala 49:25]
  assign _T_137 = _T_106[1:0]; // @[LZD.scala 49:47]
  assign _T_138 = _T_131[1:0]; // @[LZD.scala 49:59]
  assign _T_139 = _T_132 ? _T_137 : _T_138; // @[LZD.scala 49:35]
  assign _T_141 = {_T_134,_T_136,_T_139}; // @[Cat.scala 29:58]
  assign _T_142 = _T_80[3]; // @[Shift.scala 12:21]
  assign _T_143 = _T_141[3]; // @[Shift.scala 12:21]
  assign _T_144 = _T_142 | _T_143; // @[LZD.scala 49:16]
  assign _T_145 = ~ _T_143; // @[LZD.scala 49:27]
  assign _T_146 = _T_142 | _T_145; // @[LZD.scala 49:25]
  assign _T_147 = _T_80[2:0]; // @[LZD.scala 49:47]
  assign _T_148 = _T_141[2:0]; // @[LZD.scala 49:59]
  assign _T_149 = _T_142 ? _T_147 : _T_148; // @[LZD.scala 49:35]
  assign _T_151 = {_T_144,_T_146,_T_149}; // @[Cat.scala 29:58]
  assign _T_152 = _T_18[9:0]; // @[LZD.scala 44:32]
  assign _T_153 = _T_152[9:2]; // @[LZD.scala 43:32]
  assign _T_154 = _T_153[7:4]; // @[LZD.scala 43:32]
  assign _T_155 = _T_154[3:2]; // @[LZD.scala 43:32]
  assign _T_156 = _T_155 != 2'h0; // @[LZD.scala 39:14]
  assign _T_157 = _T_155[1]; // @[LZD.scala 39:21]
  assign _T_158 = _T_155[0]; // @[LZD.scala 39:30]
  assign _T_159 = ~ _T_158; // @[LZD.scala 39:27]
  assign _T_160 = _T_157 | _T_159; // @[LZD.scala 39:25]
  assign _T_161 = {_T_156,_T_160}; // @[Cat.scala 29:58]
  assign _T_162 = _T_154[1:0]; // @[LZD.scala 44:32]
  assign _T_163 = _T_162 != 2'h0; // @[LZD.scala 39:14]
  assign _T_164 = _T_162[1]; // @[LZD.scala 39:21]
  assign _T_165 = _T_162[0]; // @[LZD.scala 39:30]
  assign _T_166 = ~ _T_165; // @[LZD.scala 39:27]
  assign _T_167 = _T_164 | _T_166; // @[LZD.scala 39:25]
  assign _T_168 = {_T_163,_T_167}; // @[Cat.scala 29:58]
  assign _T_169 = _T_161[1]; // @[Shift.scala 12:21]
  assign _T_170 = _T_168[1]; // @[Shift.scala 12:21]
  assign _T_171 = _T_169 | _T_170; // @[LZD.scala 49:16]
  assign _T_172 = ~ _T_170; // @[LZD.scala 49:27]
  assign _T_173 = _T_169 | _T_172; // @[LZD.scala 49:25]
  assign _T_174 = _T_161[0:0]; // @[LZD.scala 49:47]
  assign _T_175 = _T_168[0:0]; // @[LZD.scala 49:59]
  assign _T_176 = _T_169 ? _T_174 : _T_175; // @[LZD.scala 49:35]
  assign _T_178 = {_T_171,_T_173,_T_176}; // @[Cat.scala 29:58]
  assign _T_179 = _T_153[3:0]; // @[LZD.scala 44:32]
  assign _T_180 = _T_179[3:2]; // @[LZD.scala 43:32]
  assign _T_181 = _T_180 != 2'h0; // @[LZD.scala 39:14]
  assign _T_182 = _T_180[1]; // @[LZD.scala 39:21]
  assign _T_183 = _T_180[0]; // @[LZD.scala 39:30]
  assign _T_184 = ~ _T_183; // @[LZD.scala 39:27]
  assign _T_185 = _T_182 | _T_184; // @[LZD.scala 39:25]
  assign _T_186 = {_T_181,_T_185}; // @[Cat.scala 29:58]
  assign _T_187 = _T_179[1:0]; // @[LZD.scala 44:32]
  assign _T_188 = _T_187 != 2'h0; // @[LZD.scala 39:14]
  assign _T_189 = _T_187[1]; // @[LZD.scala 39:21]
  assign _T_190 = _T_187[0]; // @[LZD.scala 39:30]
  assign _T_191 = ~ _T_190; // @[LZD.scala 39:27]
  assign _T_192 = _T_189 | _T_191; // @[LZD.scala 39:25]
  assign _T_193 = {_T_188,_T_192}; // @[Cat.scala 29:58]
  assign _T_194 = _T_186[1]; // @[Shift.scala 12:21]
  assign _T_195 = _T_193[1]; // @[Shift.scala 12:21]
  assign _T_196 = _T_194 | _T_195; // @[LZD.scala 49:16]
  assign _T_197 = ~ _T_195; // @[LZD.scala 49:27]
  assign _T_198 = _T_194 | _T_197; // @[LZD.scala 49:25]
  assign _T_199 = _T_186[0:0]; // @[LZD.scala 49:47]
  assign _T_200 = _T_193[0:0]; // @[LZD.scala 49:59]
  assign _T_201 = _T_194 ? _T_199 : _T_200; // @[LZD.scala 49:35]
  assign _T_203 = {_T_196,_T_198,_T_201}; // @[Cat.scala 29:58]
  assign _T_204 = _T_178[2]; // @[Shift.scala 12:21]
  assign _T_205 = _T_203[2]; // @[Shift.scala 12:21]
  assign _T_206 = _T_204 | _T_205; // @[LZD.scala 49:16]
  assign _T_207 = ~ _T_205; // @[LZD.scala 49:27]
  assign _T_208 = _T_204 | _T_207; // @[LZD.scala 49:25]
  assign _T_209 = _T_178[1:0]; // @[LZD.scala 49:47]
  assign _T_210 = _T_203[1:0]; // @[LZD.scala 49:59]
  assign _T_211 = _T_204 ? _T_209 : _T_210; // @[LZD.scala 49:35]
  assign _T_213 = {_T_206,_T_208,_T_211}; // @[Cat.scala 29:58]
  assign _T_214 = _T_152[1:0]; // @[LZD.scala 44:32]
  assign _T_215 = _T_214 != 2'h0; // @[LZD.scala 39:14]
  assign _T_216 = _T_214[1]; // @[LZD.scala 39:21]
  assign _T_217 = _T_214[0]; // @[LZD.scala 39:30]
  assign _T_218 = ~ _T_217; // @[LZD.scala 39:27]
  assign _T_219 = _T_216 | _T_218; // @[LZD.scala 39:25]
  assign _T_221 = _T_213[3]; // @[Shift.scala 12:21]
  assign _T_223 = {1'h1,_T_215,_T_219}; // @[Cat.scala 29:58]
  assign _T_224 = _T_213[2:0]; // @[LZD.scala 55:32]
  assign _T_225 = _T_221 ? _T_224 : _T_223; // @[LZD.scala 55:20]
  assign _T_226 = {_T_221,_T_225}; // @[Cat.scala 29:58]
  assign _T_227 = _T_151[4]; // @[Shift.scala 12:21]
  assign _T_229 = _T_151[3:0]; // @[LZD.scala 55:32]
  assign _T_230 = _T_227 ? _T_229 : _T_226; // @[LZD.scala 55:20]
  assign _T_231 = {_T_227,_T_230}; // @[Cat.scala 29:58]
  assign _T_232 = ~ _T_231; // @[convert.scala 21:22]
  assign _T_233 = realA[24:0]; // @[convert.scala 22:36]
  assign _T_234 = _T_232 < 5'h19; // @[Shift.scala 16:24]
  assign _T_236 = _T_232[4]; // @[Shift.scala 12:21]
  assign _T_237 = _T_233[8:0]; // @[Shift.scala 64:52]
  assign _T_239 = {_T_237,16'h0}; // @[Cat.scala 29:58]
  assign _T_240 = _T_236 ? _T_239 : _T_233; // @[Shift.scala 64:27]
  assign _T_241 = _T_232[3:0]; // @[Shift.scala 66:70]
  assign _T_242 = _T_241[3]; // @[Shift.scala 12:21]
  assign _T_243 = _T_240[16:0]; // @[Shift.scala 64:52]
  assign _T_245 = {_T_243,8'h0}; // @[Cat.scala 29:58]
  assign _T_246 = _T_242 ? _T_245 : _T_240; // @[Shift.scala 64:27]
  assign _T_247 = _T_241[2:0]; // @[Shift.scala 66:70]
  assign _T_248 = _T_247[2]; // @[Shift.scala 12:21]
  assign _T_249 = _T_246[20:0]; // @[Shift.scala 64:52]
  assign _T_251 = {_T_249,4'h0}; // @[Cat.scala 29:58]
  assign _T_252 = _T_248 ? _T_251 : _T_246; // @[Shift.scala 64:27]
  assign _T_253 = _T_247[1:0]; // @[Shift.scala 66:70]
  assign _T_254 = _T_253[1]; // @[Shift.scala 12:21]
  assign _T_255 = _T_252[22:0]; // @[Shift.scala 64:52]
  assign _T_257 = {_T_255,2'h0}; // @[Cat.scala 29:58]
  assign _T_258 = _T_254 ? _T_257 : _T_252; // @[Shift.scala 64:27]
  assign _T_259 = _T_253[0:0]; // @[Shift.scala 66:70]
  assign _T_261 = _T_258[23:0]; // @[Shift.scala 64:52]
  assign _T_262 = {_T_261,1'h0}; // @[Cat.scala 29:58]
  assign _T_263 = _T_259 ? _T_262 : _T_258; // @[Shift.scala 64:27]
  assign _T_264 = _T_234 ? _T_263 : 25'h0; // @[Shift.scala 16:10]
  assign _T_265 = _T_264[24:22]; // @[convert.scala 23:34]
  assign decA_fraction = _T_264[21:0]; // @[convert.scala 24:34]
  assign _T_267 = _T_15 == 1'h0; // @[convert.scala 25:26]
  assign _T_269 = _T_15 ? _T_232 : _T_231; // @[convert.scala 25:42]
  assign _T_272 = ~ _T_265; // @[convert.scala 26:67]
  assign _T_273 = _T_13 ? _T_272 : _T_265; // @[convert.scala 26:51]
  assign _T_274 = {_T_267,_T_269,_T_273}; // @[Cat.scala 29:58]
  assign _T_276 = realA[26:0]; // @[convert.scala 29:56]
  assign _T_277 = _T_276 != 27'h0; // @[convert.scala 29:60]
  assign _T_278 = ~ _T_277; // @[convert.scala 29:41]
  assign decA_isNaR = _T_13 & _T_278; // @[convert.scala 29:39]
  assign _T_281 = _T_13 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_281 & _T_278; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_274); // @[convert.scala 32:24]
  assign _T_290 = io_B[27]; // @[convert.scala 18:24]
  assign _T_291 = io_B[26]; // @[convert.scala 18:40]
  assign _T_292 = _T_290 ^ _T_291; // @[convert.scala 18:36]
  assign _T_293 = io_B[26:1]; // @[convert.scala 19:24]
  assign _T_294 = io_B[25:0]; // @[convert.scala 19:43]
  assign _T_295 = _T_293 ^ _T_294; // @[convert.scala 19:39]
  assign _T_296 = _T_295[25:10]; // @[LZD.scala 43:32]
  assign _T_297 = _T_296[15:8]; // @[LZD.scala 43:32]
  assign _T_298 = _T_297[7:4]; // @[LZD.scala 43:32]
  assign _T_299 = _T_298[3:2]; // @[LZD.scala 43:32]
  assign _T_300 = _T_299 != 2'h0; // @[LZD.scala 39:14]
  assign _T_301 = _T_299[1]; // @[LZD.scala 39:21]
  assign _T_302 = _T_299[0]; // @[LZD.scala 39:30]
  assign _T_303 = ~ _T_302; // @[LZD.scala 39:27]
  assign _T_304 = _T_301 | _T_303; // @[LZD.scala 39:25]
  assign _T_305 = {_T_300,_T_304}; // @[Cat.scala 29:58]
  assign _T_306 = _T_298[1:0]; // @[LZD.scala 44:32]
  assign _T_307 = _T_306 != 2'h0; // @[LZD.scala 39:14]
  assign _T_308 = _T_306[1]; // @[LZD.scala 39:21]
  assign _T_309 = _T_306[0]; // @[LZD.scala 39:30]
  assign _T_310 = ~ _T_309; // @[LZD.scala 39:27]
  assign _T_311 = _T_308 | _T_310; // @[LZD.scala 39:25]
  assign _T_312 = {_T_307,_T_311}; // @[Cat.scala 29:58]
  assign _T_313 = _T_305[1]; // @[Shift.scala 12:21]
  assign _T_314 = _T_312[1]; // @[Shift.scala 12:21]
  assign _T_315 = _T_313 | _T_314; // @[LZD.scala 49:16]
  assign _T_316 = ~ _T_314; // @[LZD.scala 49:27]
  assign _T_317 = _T_313 | _T_316; // @[LZD.scala 49:25]
  assign _T_318 = _T_305[0:0]; // @[LZD.scala 49:47]
  assign _T_319 = _T_312[0:0]; // @[LZD.scala 49:59]
  assign _T_320 = _T_313 ? _T_318 : _T_319; // @[LZD.scala 49:35]
  assign _T_322 = {_T_315,_T_317,_T_320}; // @[Cat.scala 29:58]
  assign _T_323 = _T_297[3:0]; // @[LZD.scala 44:32]
  assign _T_324 = _T_323[3:2]; // @[LZD.scala 43:32]
  assign _T_325 = _T_324 != 2'h0; // @[LZD.scala 39:14]
  assign _T_326 = _T_324[1]; // @[LZD.scala 39:21]
  assign _T_327 = _T_324[0]; // @[LZD.scala 39:30]
  assign _T_328 = ~ _T_327; // @[LZD.scala 39:27]
  assign _T_329 = _T_326 | _T_328; // @[LZD.scala 39:25]
  assign _T_330 = {_T_325,_T_329}; // @[Cat.scala 29:58]
  assign _T_331 = _T_323[1:0]; // @[LZD.scala 44:32]
  assign _T_332 = _T_331 != 2'h0; // @[LZD.scala 39:14]
  assign _T_333 = _T_331[1]; // @[LZD.scala 39:21]
  assign _T_334 = _T_331[0]; // @[LZD.scala 39:30]
  assign _T_335 = ~ _T_334; // @[LZD.scala 39:27]
  assign _T_336 = _T_333 | _T_335; // @[LZD.scala 39:25]
  assign _T_337 = {_T_332,_T_336}; // @[Cat.scala 29:58]
  assign _T_338 = _T_330[1]; // @[Shift.scala 12:21]
  assign _T_339 = _T_337[1]; // @[Shift.scala 12:21]
  assign _T_340 = _T_338 | _T_339; // @[LZD.scala 49:16]
  assign _T_341 = ~ _T_339; // @[LZD.scala 49:27]
  assign _T_342 = _T_338 | _T_341; // @[LZD.scala 49:25]
  assign _T_343 = _T_330[0:0]; // @[LZD.scala 49:47]
  assign _T_344 = _T_337[0:0]; // @[LZD.scala 49:59]
  assign _T_345 = _T_338 ? _T_343 : _T_344; // @[LZD.scala 49:35]
  assign _T_347 = {_T_340,_T_342,_T_345}; // @[Cat.scala 29:58]
  assign _T_348 = _T_322[2]; // @[Shift.scala 12:21]
  assign _T_349 = _T_347[2]; // @[Shift.scala 12:21]
  assign _T_350 = _T_348 | _T_349; // @[LZD.scala 49:16]
  assign _T_351 = ~ _T_349; // @[LZD.scala 49:27]
  assign _T_352 = _T_348 | _T_351; // @[LZD.scala 49:25]
  assign _T_353 = _T_322[1:0]; // @[LZD.scala 49:47]
  assign _T_354 = _T_347[1:0]; // @[LZD.scala 49:59]
  assign _T_355 = _T_348 ? _T_353 : _T_354; // @[LZD.scala 49:35]
  assign _T_357 = {_T_350,_T_352,_T_355}; // @[Cat.scala 29:58]
  assign _T_358 = _T_296[7:0]; // @[LZD.scala 44:32]
  assign _T_359 = _T_358[7:4]; // @[LZD.scala 43:32]
  assign _T_360 = _T_359[3:2]; // @[LZD.scala 43:32]
  assign _T_361 = _T_360 != 2'h0; // @[LZD.scala 39:14]
  assign _T_362 = _T_360[1]; // @[LZD.scala 39:21]
  assign _T_363 = _T_360[0]; // @[LZD.scala 39:30]
  assign _T_364 = ~ _T_363; // @[LZD.scala 39:27]
  assign _T_365 = _T_362 | _T_364; // @[LZD.scala 39:25]
  assign _T_366 = {_T_361,_T_365}; // @[Cat.scala 29:58]
  assign _T_367 = _T_359[1:0]; // @[LZD.scala 44:32]
  assign _T_368 = _T_367 != 2'h0; // @[LZD.scala 39:14]
  assign _T_369 = _T_367[1]; // @[LZD.scala 39:21]
  assign _T_370 = _T_367[0]; // @[LZD.scala 39:30]
  assign _T_371 = ~ _T_370; // @[LZD.scala 39:27]
  assign _T_372 = _T_369 | _T_371; // @[LZD.scala 39:25]
  assign _T_373 = {_T_368,_T_372}; // @[Cat.scala 29:58]
  assign _T_374 = _T_366[1]; // @[Shift.scala 12:21]
  assign _T_375 = _T_373[1]; // @[Shift.scala 12:21]
  assign _T_376 = _T_374 | _T_375; // @[LZD.scala 49:16]
  assign _T_377 = ~ _T_375; // @[LZD.scala 49:27]
  assign _T_378 = _T_374 | _T_377; // @[LZD.scala 49:25]
  assign _T_379 = _T_366[0:0]; // @[LZD.scala 49:47]
  assign _T_380 = _T_373[0:0]; // @[LZD.scala 49:59]
  assign _T_381 = _T_374 ? _T_379 : _T_380; // @[LZD.scala 49:35]
  assign _T_383 = {_T_376,_T_378,_T_381}; // @[Cat.scala 29:58]
  assign _T_384 = _T_358[3:0]; // @[LZD.scala 44:32]
  assign _T_385 = _T_384[3:2]; // @[LZD.scala 43:32]
  assign _T_386 = _T_385 != 2'h0; // @[LZD.scala 39:14]
  assign _T_387 = _T_385[1]; // @[LZD.scala 39:21]
  assign _T_388 = _T_385[0]; // @[LZD.scala 39:30]
  assign _T_389 = ~ _T_388; // @[LZD.scala 39:27]
  assign _T_390 = _T_387 | _T_389; // @[LZD.scala 39:25]
  assign _T_391 = {_T_386,_T_390}; // @[Cat.scala 29:58]
  assign _T_392 = _T_384[1:0]; // @[LZD.scala 44:32]
  assign _T_393 = _T_392 != 2'h0; // @[LZD.scala 39:14]
  assign _T_394 = _T_392[1]; // @[LZD.scala 39:21]
  assign _T_395 = _T_392[0]; // @[LZD.scala 39:30]
  assign _T_396 = ~ _T_395; // @[LZD.scala 39:27]
  assign _T_397 = _T_394 | _T_396; // @[LZD.scala 39:25]
  assign _T_398 = {_T_393,_T_397}; // @[Cat.scala 29:58]
  assign _T_399 = _T_391[1]; // @[Shift.scala 12:21]
  assign _T_400 = _T_398[1]; // @[Shift.scala 12:21]
  assign _T_401 = _T_399 | _T_400; // @[LZD.scala 49:16]
  assign _T_402 = ~ _T_400; // @[LZD.scala 49:27]
  assign _T_403 = _T_399 | _T_402; // @[LZD.scala 49:25]
  assign _T_404 = _T_391[0:0]; // @[LZD.scala 49:47]
  assign _T_405 = _T_398[0:0]; // @[LZD.scala 49:59]
  assign _T_406 = _T_399 ? _T_404 : _T_405; // @[LZD.scala 49:35]
  assign _T_408 = {_T_401,_T_403,_T_406}; // @[Cat.scala 29:58]
  assign _T_409 = _T_383[2]; // @[Shift.scala 12:21]
  assign _T_410 = _T_408[2]; // @[Shift.scala 12:21]
  assign _T_411 = _T_409 | _T_410; // @[LZD.scala 49:16]
  assign _T_412 = ~ _T_410; // @[LZD.scala 49:27]
  assign _T_413 = _T_409 | _T_412; // @[LZD.scala 49:25]
  assign _T_414 = _T_383[1:0]; // @[LZD.scala 49:47]
  assign _T_415 = _T_408[1:0]; // @[LZD.scala 49:59]
  assign _T_416 = _T_409 ? _T_414 : _T_415; // @[LZD.scala 49:35]
  assign _T_418 = {_T_411,_T_413,_T_416}; // @[Cat.scala 29:58]
  assign _T_419 = _T_357[3]; // @[Shift.scala 12:21]
  assign _T_420 = _T_418[3]; // @[Shift.scala 12:21]
  assign _T_421 = _T_419 | _T_420; // @[LZD.scala 49:16]
  assign _T_422 = ~ _T_420; // @[LZD.scala 49:27]
  assign _T_423 = _T_419 | _T_422; // @[LZD.scala 49:25]
  assign _T_424 = _T_357[2:0]; // @[LZD.scala 49:47]
  assign _T_425 = _T_418[2:0]; // @[LZD.scala 49:59]
  assign _T_426 = _T_419 ? _T_424 : _T_425; // @[LZD.scala 49:35]
  assign _T_428 = {_T_421,_T_423,_T_426}; // @[Cat.scala 29:58]
  assign _T_429 = _T_295[9:0]; // @[LZD.scala 44:32]
  assign _T_430 = _T_429[9:2]; // @[LZD.scala 43:32]
  assign _T_431 = _T_430[7:4]; // @[LZD.scala 43:32]
  assign _T_432 = _T_431[3:2]; // @[LZD.scala 43:32]
  assign _T_433 = _T_432 != 2'h0; // @[LZD.scala 39:14]
  assign _T_434 = _T_432[1]; // @[LZD.scala 39:21]
  assign _T_435 = _T_432[0]; // @[LZD.scala 39:30]
  assign _T_436 = ~ _T_435; // @[LZD.scala 39:27]
  assign _T_437 = _T_434 | _T_436; // @[LZD.scala 39:25]
  assign _T_438 = {_T_433,_T_437}; // @[Cat.scala 29:58]
  assign _T_439 = _T_431[1:0]; // @[LZD.scala 44:32]
  assign _T_440 = _T_439 != 2'h0; // @[LZD.scala 39:14]
  assign _T_441 = _T_439[1]; // @[LZD.scala 39:21]
  assign _T_442 = _T_439[0]; // @[LZD.scala 39:30]
  assign _T_443 = ~ _T_442; // @[LZD.scala 39:27]
  assign _T_444 = _T_441 | _T_443; // @[LZD.scala 39:25]
  assign _T_445 = {_T_440,_T_444}; // @[Cat.scala 29:58]
  assign _T_446 = _T_438[1]; // @[Shift.scala 12:21]
  assign _T_447 = _T_445[1]; // @[Shift.scala 12:21]
  assign _T_448 = _T_446 | _T_447; // @[LZD.scala 49:16]
  assign _T_449 = ~ _T_447; // @[LZD.scala 49:27]
  assign _T_450 = _T_446 | _T_449; // @[LZD.scala 49:25]
  assign _T_451 = _T_438[0:0]; // @[LZD.scala 49:47]
  assign _T_452 = _T_445[0:0]; // @[LZD.scala 49:59]
  assign _T_453 = _T_446 ? _T_451 : _T_452; // @[LZD.scala 49:35]
  assign _T_455 = {_T_448,_T_450,_T_453}; // @[Cat.scala 29:58]
  assign _T_456 = _T_430[3:0]; // @[LZD.scala 44:32]
  assign _T_457 = _T_456[3:2]; // @[LZD.scala 43:32]
  assign _T_458 = _T_457 != 2'h0; // @[LZD.scala 39:14]
  assign _T_459 = _T_457[1]; // @[LZD.scala 39:21]
  assign _T_460 = _T_457[0]; // @[LZD.scala 39:30]
  assign _T_461 = ~ _T_460; // @[LZD.scala 39:27]
  assign _T_462 = _T_459 | _T_461; // @[LZD.scala 39:25]
  assign _T_463 = {_T_458,_T_462}; // @[Cat.scala 29:58]
  assign _T_464 = _T_456[1:0]; // @[LZD.scala 44:32]
  assign _T_465 = _T_464 != 2'h0; // @[LZD.scala 39:14]
  assign _T_466 = _T_464[1]; // @[LZD.scala 39:21]
  assign _T_467 = _T_464[0]; // @[LZD.scala 39:30]
  assign _T_468 = ~ _T_467; // @[LZD.scala 39:27]
  assign _T_469 = _T_466 | _T_468; // @[LZD.scala 39:25]
  assign _T_470 = {_T_465,_T_469}; // @[Cat.scala 29:58]
  assign _T_471 = _T_463[1]; // @[Shift.scala 12:21]
  assign _T_472 = _T_470[1]; // @[Shift.scala 12:21]
  assign _T_473 = _T_471 | _T_472; // @[LZD.scala 49:16]
  assign _T_474 = ~ _T_472; // @[LZD.scala 49:27]
  assign _T_475 = _T_471 | _T_474; // @[LZD.scala 49:25]
  assign _T_476 = _T_463[0:0]; // @[LZD.scala 49:47]
  assign _T_477 = _T_470[0:0]; // @[LZD.scala 49:59]
  assign _T_478 = _T_471 ? _T_476 : _T_477; // @[LZD.scala 49:35]
  assign _T_480 = {_T_473,_T_475,_T_478}; // @[Cat.scala 29:58]
  assign _T_481 = _T_455[2]; // @[Shift.scala 12:21]
  assign _T_482 = _T_480[2]; // @[Shift.scala 12:21]
  assign _T_483 = _T_481 | _T_482; // @[LZD.scala 49:16]
  assign _T_484 = ~ _T_482; // @[LZD.scala 49:27]
  assign _T_485 = _T_481 | _T_484; // @[LZD.scala 49:25]
  assign _T_486 = _T_455[1:0]; // @[LZD.scala 49:47]
  assign _T_487 = _T_480[1:0]; // @[LZD.scala 49:59]
  assign _T_488 = _T_481 ? _T_486 : _T_487; // @[LZD.scala 49:35]
  assign _T_490 = {_T_483,_T_485,_T_488}; // @[Cat.scala 29:58]
  assign _T_491 = _T_429[1:0]; // @[LZD.scala 44:32]
  assign _T_492 = _T_491 != 2'h0; // @[LZD.scala 39:14]
  assign _T_493 = _T_491[1]; // @[LZD.scala 39:21]
  assign _T_494 = _T_491[0]; // @[LZD.scala 39:30]
  assign _T_495 = ~ _T_494; // @[LZD.scala 39:27]
  assign _T_496 = _T_493 | _T_495; // @[LZD.scala 39:25]
  assign _T_498 = _T_490[3]; // @[Shift.scala 12:21]
  assign _T_500 = {1'h1,_T_492,_T_496}; // @[Cat.scala 29:58]
  assign _T_501 = _T_490[2:0]; // @[LZD.scala 55:32]
  assign _T_502 = _T_498 ? _T_501 : _T_500; // @[LZD.scala 55:20]
  assign _T_503 = {_T_498,_T_502}; // @[Cat.scala 29:58]
  assign _T_504 = _T_428[4]; // @[Shift.scala 12:21]
  assign _T_506 = _T_428[3:0]; // @[LZD.scala 55:32]
  assign _T_507 = _T_504 ? _T_506 : _T_503; // @[LZD.scala 55:20]
  assign _T_508 = {_T_504,_T_507}; // @[Cat.scala 29:58]
  assign _T_509 = ~ _T_508; // @[convert.scala 21:22]
  assign _T_510 = io_B[24:0]; // @[convert.scala 22:36]
  assign _T_511 = _T_509 < 5'h19; // @[Shift.scala 16:24]
  assign _T_513 = _T_509[4]; // @[Shift.scala 12:21]
  assign _T_514 = _T_510[8:0]; // @[Shift.scala 64:52]
  assign _T_516 = {_T_514,16'h0}; // @[Cat.scala 29:58]
  assign _T_517 = _T_513 ? _T_516 : _T_510; // @[Shift.scala 64:27]
  assign _T_518 = _T_509[3:0]; // @[Shift.scala 66:70]
  assign _T_519 = _T_518[3]; // @[Shift.scala 12:21]
  assign _T_520 = _T_517[16:0]; // @[Shift.scala 64:52]
  assign _T_522 = {_T_520,8'h0}; // @[Cat.scala 29:58]
  assign _T_523 = _T_519 ? _T_522 : _T_517; // @[Shift.scala 64:27]
  assign _T_524 = _T_518[2:0]; // @[Shift.scala 66:70]
  assign _T_525 = _T_524[2]; // @[Shift.scala 12:21]
  assign _T_526 = _T_523[20:0]; // @[Shift.scala 64:52]
  assign _T_528 = {_T_526,4'h0}; // @[Cat.scala 29:58]
  assign _T_529 = _T_525 ? _T_528 : _T_523; // @[Shift.scala 64:27]
  assign _T_530 = _T_524[1:0]; // @[Shift.scala 66:70]
  assign _T_531 = _T_530[1]; // @[Shift.scala 12:21]
  assign _T_532 = _T_529[22:0]; // @[Shift.scala 64:52]
  assign _T_534 = {_T_532,2'h0}; // @[Cat.scala 29:58]
  assign _T_535 = _T_531 ? _T_534 : _T_529; // @[Shift.scala 64:27]
  assign _T_536 = _T_530[0:0]; // @[Shift.scala 66:70]
  assign _T_538 = _T_535[23:0]; // @[Shift.scala 64:52]
  assign _T_539 = {_T_538,1'h0}; // @[Cat.scala 29:58]
  assign _T_540 = _T_536 ? _T_539 : _T_535; // @[Shift.scala 64:27]
  assign _T_541 = _T_511 ? _T_540 : 25'h0; // @[Shift.scala 16:10]
  assign _T_542 = _T_541[24:22]; // @[convert.scala 23:34]
  assign decB_fraction = _T_541[21:0]; // @[convert.scala 24:34]
  assign _T_544 = _T_292 == 1'h0; // @[convert.scala 25:26]
  assign _T_546 = _T_292 ? _T_509 : _T_508; // @[convert.scala 25:42]
  assign _T_549 = ~ _T_542; // @[convert.scala 26:67]
  assign _T_550 = _T_290 ? _T_549 : _T_542; // @[convert.scala 26:51]
  assign _T_551 = {_T_544,_T_546,_T_550}; // @[Cat.scala 29:58]
  assign _T_553 = io_B[26:0]; // @[convert.scala 29:56]
  assign _T_554 = _T_553 != 27'h0; // @[convert.scala 29:60]
  assign _T_555 = ~ _T_554; // @[convert.scala 29:41]
  assign decB_isNaR = _T_290 & _T_555; // @[convert.scala 29:39]
  assign _T_558 = _T_290 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_558 & _T_555; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_551); // @[convert.scala 32:24]
  assign _T_567 = realC[27]; // @[convert.scala 18:24]
  assign _T_568 = realC[26]; // @[convert.scala 18:40]
  assign _T_569 = _T_567 ^ _T_568; // @[convert.scala 18:36]
  assign _T_570 = realC[26:1]; // @[convert.scala 19:24]
  assign _T_571 = realC[25:0]; // @[convert.scala 19:43]
  assign _T_572 = _T_570 ^ _T_571; // @[convert.scala 19:39]
  assign _T_573 = _T_572[25:10]; // @[LZD.scala 43:32]
  assign _T_574 = _T_573[15:8]; // @[LZD.scala 43:32]
  assign _T_575 = _T_574[7:4]; // @[LZD.scala 43:32]
  assign _T_576 = _T_575[3:2]; // @[LZD.scala 43:32]
  assign _T_577 = _T_576 != 2'h0; // @[LZD.scala 39:14]
  assign _T_578 = _T_576[1]; // @[LZD.scala 39:21]
  assign _T_579 = _T_576[0]; // @[LZD.scala 39:30]
  assign _T_580 = ~ _T_579; // @[LZD.scala 39:27]
  assign _T_581 = _T_578 | _T_580; // @[LZD.scala 39:25]
  assign _T_582 = {_T_577,_T_581}; // @[Cat.scala 29:58]
  assign _T_583 = _T_575[1:0]; // @[LZD.scala 44:32]
  assign _T_584 = _T_583 != 2'h0; // @[LZD.scala 39:14]
  assign _T_585 = _T_583[1]; // @[LZD.scala 39:21]
  assign _T_586 = _T_583[0]; // @[LZD.scala 39:30]
  assign _T_587 = ~ _T_586; // @[LZD.scala 39:27]
  assign _T_588 = _T_585 | _T_587; // @[LZD.scala 39:25]
  assign _T_589 = {_T_584,_T_588}; // @[Cat.scala 29:58]
  assign _T_590 = _T_582[1]; // @[Shift.scala 12:21]
  assign _T_591 = _T_589[1]; // @[Shift.scala 12:21]
  assign _T_592 = _T_590 | _T_591; // @[LZD.scala 49:16]
  assign _T_593 = ~ _T_591; // @[LZD.scala 49:27]
  assign _T_594 = _T_590 | _T_593; // @[LZD.scala 49:25]
  assign _T_595 = _T_582[0:0]; // @[LZD.scala 49:47]
  assign _T_596 = _T_589[0:0]; // @[LZD.scala 49:59]
  assign _T_597 = _T_590 ? _T_595 : _T_596; // @[LZD.scala 49:35]
  assign _T_599 = {_T_592,_T_594,_T_597}; // @[Cat.scala 29:58]
  assign _T_600 = _T_574[3:0]; // @[LZD.scala 44:32]
  assign _T_601 = _T_600[3:2]; // @[LZD.scala 43:32]
  assign _T_602 = _T_601 != 2'h0; // @[LZD.scala 39:14]
  assign _T_603 = _T_601[1]; // @[LZD.scala 39:21]
  assign _T_604 = _T_601[0]; // @[LZD.scala 39:30]
  assign _T_605 = ~ _T_604; // @[LZD.scala 39:27]
  assign _T_606 = _T_603 | _T_605; // @[LZD.scala 39:25]
  assign _T_607 = {_T_602,_T_606}; // @[Cat.scala 29:58]
  assign _T_608 = _T_600[1:0]; // @[LZD.scala 44:32]
  assign _T_609 = _T_608 != 2'h0; // @[LZD.scala 39:14]
  assign _T_610 = _T_608[1]; // @[LZD.scala 39:21]
  assign _T_611 = _T_608[0]; // @[LZD.scala 39:30]
  assign _T_612 = ~ _T_611; // @[LZD.scala 39:27]
  assign _T_613 = _T_610 | _T_612; // @[LZD.scala 39:25]
  assign _T_614 = {_T_609,_T_613}; // @[Cat.scala 29:58]
  assign _T_615 = _T_607[1]; // @[Shift.scala 12:21]
  assign _T_616 = _T_614[1]; // @[Shift.scala 12:21]
  assign _T_617 = _T_615 | _T_616; // @[LZD.scala 49:16]
  assign _T_618 = ~ _T_616; // @[LZD.scala 49:27]
  assign _T_619 = _T_615 | _T_618; // @[LZD.scala 49:25]
  assign _T_620 = _T_607[0:0]; // @[LZD.scala 49:47]
  assign _T_621 = _T_614[0:0]; // @[LZD.scala 49:59]
  assign _T_622 = _T_615 ? _T_620 : _T_621; // @[LZD.scala 49:35]
  assign _T_624 = {_T_617,_T_619,_T_622}; // @[Cat.scala 29:58]
  assign _T_625 = _T_599[2]; // @[Shift.scala 12:21]
  assign _T_626 = _T_624[2]; // @[Shift.scala 12:21]
  assign _T_627 = _T_625 | _T_626; // @[LZD.scala 49:16]
  assign _T_628 = ~ _T_626; // @[LZD.scala 49:27]
  assign _T_629 = _T_625 | _T_628; // @[LZD.scala 49:25]
  assign _T_630 = _T_599[1:0]; // @[LZD.scala 49:47]
  assign _T_631 = _T_624[1:0]; // @[LZD.scala 49:59]
  assign _T_632 = _T_625 ? _T_630 : _T_631; // @[LZD.scala 49:35]
  assign _T_634 = {_T_627,_T_629,_T_632}; // @[Cat.scala 29:58]
  assign _T_635 = _T_573[7:0]; // @[LZD.scala 44:32]
  assign _T_636 = _T_635[7:4]; // @[LZD.scala 43:32]
  assign _T_637 = _T_636[3:2]; // @[LZD.scala 43:32]
  assign _T_638 = _T_637 != 2'h0; // @[LZD.scala 39:14]
  assign _T_639 = _T_637[1]; // @[LZD.scala 39:21]
  assign _T_640 = _T_637[0]; // @[LZD.scala 39:30]
  assign _T_641 = ~ _T_640; // @[LZD.scala 39:27]
  assign _T_642 = _T_639 | _T_641; // @[LZD.scala 39:25]
  assign _T_643 = {_T_638,_T_642}; // @[Cat.scala 29:58]
  assign _T_644 = _T_636[1:0]; // @[LZD.scala 44:32]
  assign _T_645 = _T_644 != 2'h0; // @[LZD.scala 39:14]
  assign _T_646 = _T_644[1]; // @[LZD.scala 39:21]
  assign _T_647 = _T_644[0]; // @[LZD.scala 39:30]
  assign _T_648 = ~ _T_647; // @[LZD.scala 39:27]
  assign _T_649 = _T_646 | _T_648; // @[LZD.scala 39:25]
  assign _T_650 = {_T_645,_T_649}; // @[Cat.scala 29:58]
  assign _T_651 = _T_643[1]; // @[Shift.scala 12:21]
  assign _T_652 = _T_650[1]; // @[Shift.scala 12:21]
  assign _T_653 = _T_651 | _T_652; // @[LZD.scala 49:16]
  assign _T_654 = ~ _T_652; // @[LZD.scala 49:27]
  assign _T_655 = _T_651 | _T_654; // @[LZD.scala 49:25]
  assign _T_656 = _T_643[0:0]; // @[LZD.scala 49:47]
  assign _T_657 = _T_650[0:0]; // @[LZD.scala 49:59]
  assign _T_658 = _T_651 ? _T_656 : _T_657; // @[LZD.scala 49:35]
  assign _T_660 = {_T_653,_T_655,_T_658}; // @[Cat.scala 29:58]
  assign _T_661 = _T_635[3:0]; // @[LZD.scala 44:32]
  assign _T_662 = _T_661[3:2]; // @[LZD.scala 43:32]
  assign _T_663 = _T_662 != 2'h0; // @[LZD.scala 39:14]
  assign _T_664 = _T_662[1]; // @[LZD.scala 39:21]
  assign _T_665 = _T_662[0]; // @[LZD.scala 39:30]
  assign _T_666 = ~ _T_665; // @[LZD.scala 39:27]
  assign _T_667 = _T_664 | _T_666; // @[LZD.scala 39:25]
  assign _T_668 = {_T_663,_T_667}; // @[Cat.scala 29:58]
  assign _T_669 = _T_661[1:0]; // @[LZD.scala 44:32]
  assign _T_670 = _T_669 != 2'h0; // @[LZD.scala 39:14]
  assign _T_671 = _T_669[1]; // @[LZD.scala 39:21]
  assign _T_672 = _T_669[0]; // @[LZD.scala 39:30]
  assign _T_673 = ~ _T_672; // @[LZD.scala 39:27]
  assign _T_674 = _T_671 | _T_673; // @[LZD.scala 39:25]
  assign _T_675 = {_T_670,_T_674}; // @[Cat.scala 29:58]
  assign _T_676 = _T_668[1]; // @[Shift.scala 12:21]
  assign _T_677 = _T_675[1]; // @[Shift.scala 12:21]
  assign _T_678 = _T_676 | _T_677; // @[LZD.scala 49:16]
  assign _T_679 = ~ _T_677; // @[LZD.scala 49:27]
  assign _T_680 = _T_676 | _T_679; // @[LZD.scala 49:25]
  assign _T_681 = _T_668[0:0]; // @[LZD.scala 49:47]
  assign _T_682 = _T_675[0:0]; // @[LZD.scala 49:59]
  assign _T_683 = _T_676 ? _T_681 : _T_682; // @[LZD.scala 49:35]
  assign _T_685 = {_T_678,_T_680,_T_683}; // @[Cat.scala 29:58]
  assign _T_686 = _T_660[2]; // @[Shift.scala 12:21]
  assign _T_687 = _T_685[2]; // @[Shift.scala 12:21]
  assign _T_688 = _T_686 | _T_687; // @[LZD.scala 49:16]
  assign _T_689 = ~ _T_687; // @[LZD.scala 49:27]
  assign _T_690 = _T_686 | _T_689; // @[LZD.scala 49:25]
  assign _T_691 = _T_660[1:0]; // @[LZD.scala 49:47]
  assign _T_692 = _T_685[1:0]; // @[LZD.scala 49:59]
  assign _T_693 = _T_686 ? _T_691 : _T_692; // @[LZD.scala 49:35]
  assign _T_695 = {_T_688,_T_690,_T_693}; // @[Cat.scala 29:58]
  assign _T_696 = _T_634[3]; // @[Shift.scala 12:21]
  assign _T_697 = _T_695[3]; // @[Shift.scala 12:21]
  assign _T_698 = _T_696 | _T_697; // @[LZD.scala 49:16]
  assign _T_699 = ~ _T_697; // @[LZD.scala 49:27]
  assign _T_700 = _T_696 | _T_699; // @[LZD.scala 49:25]
  assign _T_701 = _T_634[2:0]; // @[LZD.scala 49:47]
  assign _T_702 = _T_695[2:0]; // @[LZD.scala 49:59]
  assign _T_703 = _T_696 ? _T_701 : _T_702; // @[LZD.scala 49:35]
  assign _T_705 = {_T_698,_T_700,_T_703}; // @[Cat.scala 29:58]
  assign _T_706 = _T_572[9:0]; // @[LZD.scala 44:32]
  assign _T_707 = _T_706[9:2]; // @[LZD.scala 43:32]
  assign _T_708 = _T_707[7:4]; // @[LZD.scala 43:32]
  assign _T_709 = _T_708[3:2]; // @[LZD.scala 43:32]
  assign _T_710 = _T_709 != 2'h0; // @[LZD.scala 39:14]
  assign _T_711 = _T_709[1]; // @[LZD.scala 39:21]
  assign _T_712 = _T_709[0]; // @[LZD.scala 39:30]
  assign _T_713 = ~ _T_712; // @[LZD.scala 39:27]
  assign _T_714 = _T_711 | _T_713; // @[LZD.scala 39:25]
  assign _T_715 = {_T_710,_T_714}; // @[Cat.scala 29:58]
  assign _T_716 = _T_708[1:0]; // @[LZD.scala 44:32]
  assign _T_717 = _T_716 != 2'h0; // @[LZD.scala 39:14]
  assign _T_718 = _T_716[1]; // @[LZD.scala 39:21]
  assign _T_719 = _T_716[0]; // @[LZD.scala 39:30]
  assign _T_720 = ~ _T_719; // @[LZD.scala 39:27]
  assign _T_721 = _T_718 | _T_720; // @[LZD.scala 39:25]
  assign _T_722 = {_T_717,_T_721}; // @[Cat.scala 29:58]
  assign _T_723 = _T_715[1]; // @[Shift.scala 12:21]
  assign _T_724 = _T_722[1]; // @[Shift.scala 12:21]
  assign _T_725 = _T_723 | _T_724; // @[LZD.scala 49:16]
  assign _T_726 = ~ _T_724; // @[LZD.scala 49:27]
  assign _T_727 = _T_723 | _T_726; // @[LZD.scala 49:25]
  assign _T_728 = _T_715[0:0]; // @[LZD.scala 49:47]
  assign _T_729 = _T_722[0:0]; // @[LZD.scala 49:59]
  assign _T_730 = _T_723 ? _T_728 : _T_729; // @[LZD.scala 49:35]
  assign _T_732 = {_T_725,_T_727,_T_730}; // @[Cat.scala 29:58]
  assign _T_733 = _T_707[3:0]; // @[LZD.scala 44:32]
  assign _T_734 = _T_733[3:2]; // @[LZD.scala 43:32]
  assign _T_735 = _T_734 != 2'h0; // @[LZD.scala 39:14]
  assign _T_736 = _T_734[1]; // @[LZD.scala 39:21]
  assign _T_737 = _T_734[0]; // @[LZD.scala 39:30]
  assign _T_738 = ~ _T_737; // @[LZD.scala 39:27]
  assign _T_739 = _T_736 | _T_738; // @[LZD.scala 39:25]
  assign _T_740 = {_T_735,_T_739}; // @[Cat.scala 29:58]
  assign _T_741 = _T_733[1:0]; // @[LZD.scala 44:32]
  assign _T_742 = _T_741 != 2'h0; // @[LZD.scala 39:14]
  assign _T_743 = _T_741[1]; // @[LZD.scala 39:21]
  assign _T_744 = _T_741[0]; // @[LZD.scala 39:30]
  assign _T_745 = ~ _T_744; // @[LZD.scala 39:27]
  assign _T_746 = _T_743 | _T_745; // @[LZD.scala 39:25]
  assign _T_747 = {_T_742,_T_746}; // @[Cat.scala 29:58]
  assign _T_748 = _T_740[1]; // @[Shift.scala 12:21]
  assign _T_749 = _T_747[1]; // @[Shift.scala 12:21]
  assign _T_750 = _T_748 | _T_749; // @[LZD.scala 49:16]
  assign _T_751 = ~ _T_749; // @[LZD.scala 49:27]
  assign _T_752 = _T_748 | _T_751; // @[LZD.scala 49:25]
  assign _T_753 = _T_740[0:0]; // @[LZD.scala 49:47]
  assign _T_754 = _T_747[0:0]; // @[LZD.scala 49:59]
  assign _T_755 = _T_748 ? _T_753 : _T_754; // @[LZD.scala 49:35]
  assign _T_757 = {_T_750,_T_752,_T_755}; // @[Cat.scala 29:58]
  assign _T_758 = _T_732[2]; // @[Shift.scala 12:21]
  assign _T_759 = _T_757[2]; // @[Shift.scala 12:21]
  assign _T_760 = _T_758 | _T_759; // @[LZD.scala 49:16]
  assign _T_761 = ~ _T_759; // @[LZD.scala 49:27]
  assign _T_762 = _T_758 | _T_761; // @[LZD.scala 49:25]
  assign _T_763 = _T_732[1:0]; // @[LZD.scala 49:47]
  assign _T_764 = _T_757[1:0]; // @[LZD.scala 49:59]
  assign _T_765 = _T_758 ? _T_763 : _T_764; // @[LZD.scala 49:35]
  assign _T_767 = {_T_760,_T_762,_T_765}; // @[Cat.scala 29:58]
  assign _T_768 = _T_706[1:0]; // @[LZD.scala 44:32]
  assign _T_769 = _T_768 != 2'h0; // @[LZD.scala 39:14]
  assign _T_770 = _T_768[1]; // @[LZD.scala 39:21]
  assign _T_771 = _T_768[0]; // @[LZD.scala 39:30]
  assign _T_772 = ~ _T_771; // @[LZD.scala 39:27]
  assign _T_773 = _T_770 | _T_772; // @[LZD.scala 39:25]
  assign _T_775 = _T_767[3]; // @[Shift.scala 12:21]
  assign _T_777 = {1'h1,_T_769,_T_773}; // @[Cat.scala 29:58]
  assign _T_778 = _T_767[2:0]; // @[LZD.scala 55:32]
  assign _T_779 = _T_775 ? _T_778 : _T_777; // @[LZD.scala 55:20]
  assign _T_780 = {_T_775,_T_779}; // @[Cat.scala 29:58]
  assign _T_781 = _T_705[4]; // @[Shift.scala 12:21]
  assign _T_783 = _T_705[3:0]; // @[LZD.scala 55:32]
  assign _T_784 = _T_781 ? _T_783 : _T_780; // @[LZD.scala 55:20]
  assign _T_785 = {_T_781,_T_784}; // @[Cat.scala 29:58]
  assign _T_786 = ~ _T_785; // @[convert.scala 21:22]
  assign _T_787 = realC[24:0]; // @[convert.scala 22:36]
  assign _T_788 = _T_786 < 5'h19; // @[Shift.scala 16:24]
  assign _T_790 = _T_786[4]; // @[Shift.scala 12:21]
  assign _T_791 = _T_787[8:0]; // @[Shift.scala 64:52]
  assign _T_793 = {_T_791,16'h0}; // @[Cat.scala 29:58]
  assign _T_794 = _T_790 ? _T_793 : _T_787; // @[Shift.scala 64:27]
  assign _T_795 = _T_786[3:0]; // @[Shift.scala 66:70]
  assign _T_796 = _T_795[3]; // @[Shift.scala 12:21]
  assign _T_797 = _T_794[16:0]; // @[Shift.scala 64:52]
  assign _T_799 = {_T_797,8'h0}; // @[Cat.scala 29:58]
  assign _T_800 = _T_796 ? _T_799 : _T_794; // @[Shift.scala 64:27]
  assign _T_801 = _T_795[2:0]; // @[Shift.scala 66:70]
  assign _T_802 = _T_801[2]; // @[Shift.scala 12:21]
  assign _T_803 = _T_800[20:0]; // @[Shift.scala 64:52]
  assign _T_805 = {_T_803,4'h0}; // @[Cat.scala 29:58]
  assign _T_806 = _T_802 ? _T_805 : _T_800; // @[Shift.scala 64:27]
  assign _T_807 = _T_801[1:0]; // @[Shift.scala 66:70]
  assign _T_808 = _T_807[1]; // @[Shift.scala 12:21]
  assign _T_809 = _T_806[22:0]; // @[Shift.scala 64:52]
  assign _T_811 = {_T_809,2'h0}; // @[Cat.scala 29:58]
  assign _T_812 = _T_808 ? _T_811 : _T_806; // @[Shift.scala 64:27]
  assign _T_813 = _T_807[0:0]; // @[Shift.scala 66:70]
  assign _T_815 = _T_812[23:0]; // @[Shift.scala 64:52]
  assign _T_816 = {_T_815,1'h0}; // @[Cat.scala 29:58]
  assign _T_817 = _T_813 ? _T_816 : _T_812; // @[Shift.scala 64:27]
  assign _T_818 = _T_788 ? _T_817 : 25'h0; // @[Shift.scala 16:10]
  assign _T_819 = _T_818[24:22]; // @[convert.scala 23:34]
  assign decC_fraction = _T_818[21:0]; // @[convert.scala 24:34]
  assign _T_821 = _T_569 == 1'h0; // @[convert.scala 25:26]
  assign _T_823 = _T_569 ? _T_786 : _T_785; // @[convert.scala 25:42]
  assign _T_826 = ~ _T_819; // @[convert.scala 26:67]
  assign _T_827 = _T_567 ? _T_826 : _T_819; // @[convert.scala 26:51]
  assign _T_828 = {_T_821,_T_823,_T_827}; // @[Cat.scala 29:58]
  assign _T_830 = realC[26:0]; // @[convert.scala 29:56]
  assign _T_831 = _T_830 != 27'h0; // @[convert.scala 29:60]
  assign _T_832 = ~ _T_831; // @[convert.scala 29:41]
  assign decC_isNaR = _T_567 & _T_832; // @[convert.scala 29:39]
  assign _T_835 = _T_567 == 1'h0; // @[convert.scala 30:19]
  assign decC_isZero = _T_835 & _T_832; // @[convert.scala 30:41]
  assign decC_scale = $signed(_T_828); // @[convert.scala 32:24]
  assign _T_843 = decA_isNaR | decB_isNaR; // @[PositFMA.scala 58:30]
  assign outIsNaR = _T_843 | decC_isNaR; // @[PositFMA.scala 58:44]
  assign _T_844 = ~ _T_13; // @[PositFMA.scala 59:34]
  assign _T_845 = ~ decA_isZero; // @[PositFMA.scala 59:47]
  assign _T_846 = _T_844 & _T_845; // @[PositFMA.scala 59:45]
  assign _T_848 = {_T_13,_T_846,decA_fraction}; // @[Cat.scala 29:58]
  assign sigA = $signed(_T_848); // @[PositFMA.scala 59:76]
  assign _T_849 = ~ _T_290; // @[PositFMA.scala 60:34]
  assign _T_850 = ~ decB_isZero; // @[PositFMA.scala 60:47]
  assign _T_851 = _T_849 & _T_850; // @[PositFMA.scala 60:45]
  assign _T_853 = {_T_290,_T_851,decB_fraction}; // @[Cat.scala 29:58]
  assign sigB = $signed(_T_853); // @[PositFMA.scala 60:76]
  assign _T_854 = $signed(sigA) * $signed(sigB); // @[PositFMA.scala 61:25]
  assign sigP = $unsigned(_T_854); // @[PositFMA.scala 61:33]
  assign head2 = sigP[47:46]; // @[PositFMA.scala 62:28]
  assign _T_855 = head2[1]; // @[PositFMA.scala 63:31]
  assign _T_856 = ~ _T_855; // @[PositFMA.scala 63:25]
  assign _T_857 = head2[0]; // @[PositFMA.scala 63:42]
  assign addTwo = _T_856 & _T_857; // @[PositFMA.scala 63:35]
  assign _T_858 = sigP[47]; // @[PositFMA.scala 65:23]
  assign _T_859 = sigP[45]; // @[PositFMA.scala 65:49]
  assign addOne = _T_858 ^ _T_859; // @[PositFMA.scala 65:43]
  assign _T_860 = {addTwo,addOne}; // @[Cat.scala 29:58]
  assign expBias = {1'b0,$signed(_T_860)}; // @[PositFMA.scala 66:39]
  assign mulSign = sigP[47:47]; // @[PositFMA.scala 67:28]
  assign _T_861 = $signed(decA_scale) + $signed(decB_scale); // @[PositFMA.scala 69:30]
  assign _GEN_12 = {{7{expBias[2]}},expBias}; // @[PositFMA.scala 69:44]
  assign _T_863 = $signed(_T_861) + $signed(_GEN_12); // @[PositFMA.scala 69:44]
  assign mulScale = $signed(_T_863); // @[PositFMA.scala 69:44]
  assign _T_864 = sigP[45:0]; // @[PositFMA.scala 72:29]
  assign _T_865 = sigP[44:0]; // @[PositFMA.scala 73:29]
  assign _T_866 = {_T_865, 1'h0}; // @[PositFMA.scala 73:48]
  assign mulSigTmp = addOne ? _T_864 : _T_866; // @[PositFMA.scala 70:22]
  assign _T_868 = mulSigTmp[45:45]; // @[PositFMA.scala 77:39]
  assign _T_869 = _T_868 | addTwo; // @[PositFMA.scala 77:43]
  assign _T_870 = mulSigTmp[44:0]; // @[PositFMA.scala 78:39]
  assign mulSig = {mulSign,_T_869,_T_870}; // @[Cat.scala 29:58]
  assign _T_896 = ~ addSign_phase2; // @[PositFMA.scala 107:29]
  assign _T_897 = ~ addZero_phase2; // @[PositFMA.scala 107:47]
  assign _T_898 = _T_896 & _T_897; // @[PositFMA.scala 107:45]
  assign extAddSig = {addSign_phase2,_T_898,addFrac_phase2,23'h0}; // @[Cat.scala 29:58]
  assign _GEN_13 = {{1{addScale_phase2[8]}},addScale_phase2}; // @[PositFMA.scala 111:39]
  assign mulGreater = $signed(mulScale_phase2) > $signed(_GEN_13); // @[PositFMA.scala 111:39]
  assign greaterScale = mulGreater ? $signed(mulScale_phase2) : $signed({{1{addScale_phase2[8]}},addScale_phase2}); // @[PositFMA.scala 112:26]
  assign smallerScale = mulGreater ? $signed({{1{addScale_phase2[8]}},addScale_phase2}) : $signed(mulScale_phase2); // @[PositFMA.scala 113:26]
  assign _T_902 = $signed(greaterScale) - $signed(smallerScale); // @[PositFMA.scala 114:36]
  assign scaleDiff = $signed(_T_902); // @[PositFMA.scala 114:36]
  assign greaterSig = mulGreater ? mulSig_phase2 : extAddSig; // @[PositFMA.scala 115:26]
  assign smallerSigTmp = mulGreater ? extAddSig : mulSig_phase2; // @[PositFMA.scala 116:26]
  assign _T_903 = $unsigned(scaleDiff); // @[PositFMA.scala 117:69]
  assign _T_904 = _T_903 < 10'h2f; // @[Shift.scala 39:24]
  assign _T_905 = _T_903[5:0]; // @[Shift.scala 40:44]
  assign _T_906 = smallerSigTmp[46:32]; // @[Shift.scala 90:30]
  assign _T_907 = smallerSigTmp[31:0]; // @[Shift.scala 90:48]
  assign _T_908 = _T_907 != 32'h0; // @[Shift.scala 90:57]
  assign _GEN_14 = {{14'd0}, _T_908}; // @[Shift.scala 90:39]
  assign _T_909 = _T_906 | _GEN_14; // @[Shift.scala 90:39]
  assign _T_910 = _T_905[5]; // @[Shift.scala 12:21]
  assign _T_911 = smallerSigTmp[46]; // @[Shift.scala 12:21]
  assign _T_913 = _T_911 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 71:12]
  assign _T_914 = {_T_913,_T_909}; // @[Cat.scala 29:58]
  assign _T_915 = _T_910 ? _T_914 : smallerSigTmp; // @[Shift.scala 91:22]
  assign _T_916 = _T_905[4:0]; // @[Shift.scala 92:77]
  assign _T_917 = _T_915[46:16]; // @[Shift.scala 90:30]
  assign _T_918 = _T_915[15:0]; // @[Shift.scala 90:48]
  assign _T_919 = _T_918 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_15 = {{30'd0}, _T_919}; // @[Shift.scala 90:39]
  assign _T_920 = _T_917 | _GEN_15; // @[Shift.scala 90:39]
  assign _T_921 = _T_916[4]; // @[Shift.scala 12:21]
  assign _T_922 = _T_915[46]; // @[Shift.scala 12:21]
  assign _T_924 = _T_922 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_925 = {_T_924,_T_920}; // @[Cat.scala 29:58]
  assign _T_926 = _T_921 ? _T_925 : _T_915; // @[Shift.scala 91:22]
  assign _T_927 = _T_916[3:0]; // @[Shift.scala 92:77]
  assign _T_928 = _T_926[46:8]; // @[Shift.scala 90:30]
  assign _T_929 = _T_926[7:0]; // @[Shift.scala 90:48]
  assign _T_930 = _T_929 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_16 = {{38'd0}, _T_930}; // @[Shift.scala 90:39]
  assign _T_931 = _T_928 | _GEN_16; // @[Shift.scala 90:39]
  assign _T_932 = _T_927[3]; // @[Shift.scala 12:21]
  assign _T_933 = _T_926[46]; // @[Shift.scala 12:21]
  assign _T_935 = _T_933 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_936 = {_T_935,_T_931}; // @[Cat.scala 29:58]
  assign _T_937 = _T_932 ? _T_936 : _T_926; // @[Shift.scala 91:22]
  assign _T_938 = _T_927[2:0]; // @[Shift.scala 92:77]
  assign _T_939 = _T_937[46:4]; // @[Shift.scala 90:30]
  assign _T_940 = _T_937[3:0]; // @[Shift.scala 90:48]
  assign _T_941 = _T_940 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_17 = {{42'd0}, _T_941}; // @[Shift.scala 90:39]
  assign _T_942 = _T_939 | _GEN_17; // @[Shift.scala 90:39]
  assign _T_943 = _T_938[2]; // @[Shift.scala 12:21]
  assign _T_944 = _T_937[46]; // @[Shift.scala 12:21]
  assign _T_946 = _T_944 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_947 = {_T_946,_T_942}; // @[Cat.scala 29:58]
  assign _T_948 = _T_943 ? _T_947 : _T_937; // @[Shift.scala 91:22]
  assign _T_949 = _T_938[1:0]; // @[Shift.scala 92:77]
  assign _T_950 = _T_948[46:2]; // @[Shift.scala 90:30]
  assign _T_951 = _T_948[1:0]; // @[Shift.scala 90:48]
  assign _T_952 = _T_951 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_18 = {{44'd0}, _T_952}; // @[Shift.scala 90:39]
  assign _T_953 = _T_950 | _GEN_18; // @[Shift.scala 90:39]
  assign _T_954 = _T_949[1]; // @[Shift.scala 12:21]
  assign _T_955 = _T_948[46]; // @[Shift.scala 12:21]
  assign _T_957 = _T_955 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_958 = {_T_957,_T_953}; // @[Cat.scala 29:58]
  assign _T_959 = _T_954 ? _T_958 : _T_948; // @[Shift.scala 91:22]
  assign _T_960 = _T_949[0:0]; // @[Shift.scala 92:77]
  assign _T_961 = _T_959[46:1]; // @[Shift.scala 90:30]
  assign _T_962 = _T_959[0:0]; // @[Shift.scala 90:48]
  assign _GEN_19 = {{45'd0}, _T_962}; // @[Shift.scala 90:39]
  assign _T_964 = _T_961 | _GEN_19; // @[Shift.scala 90:39]
  assign _T_966 = _T_959[46]; // @[Shift.scala 12:21]
  assign _T_967 = {_T_966,_T_964}; // @[Cat.scala 29:58]
  assign _T_968 = _T_960 ? _T_967 : _T_959; // @[Shift.scala 91:22]
  assign _T_971 = _T_911 ? 47'h7fffffffffff : 47'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_904 ? _T_968 : _T_971; // @[Shift.scala 39:10]
  assign rawSumSig = greaterSig + smallerSig; // @[PositFMA.scala 118:34]
  assign _T_972 = mulSig_phase2[46:46]; // @[PositFMA.scala 119:42]
  assign _T_973 = _T_972 ^ addSign_phase2; // @[PositFMA.scala 119:46]
  assign _T_974 = rawSumSig[47:47]; // @[PositFMA.scala 119:79]
  assign sumSign = _T_973 ^ _T_974; // @[PositFMA.scala 119:63]
  assign _T_976 = greaterSig + smallerSig; // @[PositFMA.scala 120:50]
  assign signSumSig = {sumSign,_T_976}; // @[Cat.scala 29:58]
  assign _T_977 = signSumSig[47:1]; // @[PositFMA.scala 124:33]
  assign _T_978 = signSumSig[46:0]; // @[PositFMA.scala 124:68]
  assign sumXor = _T_977 ^ _T_978; // @[PositFMA.scala 124:51]
  assign _T_979 = sumXor[46:15]; // @[LZD.scala 43:32]
  assign _T_980 = _T_979[31:16]; // @[LZD.scala 43:32]
  assign _T_981 = _T_980[15:8]; // @[LZD.scala 43:32]
  assign _T_982 = _T_981[7:4]; // @[LZD.scala 43:32]
  assign _T_983 = _T_982[3:2]; // @[LZD.scala 43:32]
  assign _T_984 = _T_983 != 2'h0; // @[LZD.scala 39:14]
  assign _T_985 = _T_983[1]; // @[LZD.scala 39:21]
  assign _T_986 = _T_983[0]; // @[LZD.scala 39:30]
  assign _T_987 = ~ _T_986; // @[LZD.scala 39:27]
  assign _T_988 = _T_985 | _T_987; // @[LZD.scala 39:25]
  assign _T_989 = {_T_984,_T_988}; // @[Cat.scala 29:58]
  assign _T_990 = _T_982[1:0]; // @[LZD.scala 44:32]
  assign _T_991 = _T_990 != 2'h0; // @[LZD.scala 39:14]
  assign _T_992 = _T_990[1]; // @[LZD.scala 39:21]
  assign _T_993 = _T_990[0]; // @[LZD.scala 39:30]
  assign _T_994 = ~ _T_993; // @[LZD.scala 39:27]
  assign _T_995 = _T_992 | _T_994; // @[LZD.scala 39:25]
  assign _T_996 = {_T_991,_T_995}; // @[Cat.scala 29:58]
  assign _T_997 = _T_989[1]; // @[Shift.scala 12:21]
  assign _T_998 = _T_996[1]; // @[Shift.scala 12:21]
  assign _T_999 = _T_997 | _T_998; // @[LZD.scala 49:16]
  assign _T_1000 = ~ _T_998; // @[LZD.scala 49:27]
  assign _T_1001 = _T_997 | _T_1000; // @[LZD.scala 49:25]
  assign _T_1002 = _T_989[0:0]; // @[LZD.scala 49:47]
  assign _T_1003 = _T_996[0:0]; // @[LZD.scala 49:59]
  assign _T_1004 = _T_997 ? _T_1002 : _T_1003; // @[LZD.scala 49:35]
  assign _T_1006 = {_T_999,_T_1001,_T_1004}; // @[Cat.scala 29:58]
  assign _T_1007 = _T_981[3:0]; // @[LZD.scala 44:32]
  assign _T_1008 = _T_1007[3:2]; // @[LZD.scala 43:32]
  assign _T_1009 = _T_1008 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1010 = _T_1008[1]; // @[LZD.scala 39:21]
  assign _T_1011 = _T_1008[0]; // @[LZD.scala 39:30]
  assign _T_1012 = ~ _T_1011; // @[LZD.scala 39:27]
  assign _T_1013 = _T_1010 | _T_1012; // @[LZD.scala 39:25]
  assign _T_1014 = {_T_1009,_T_1013}; // @[Cat.scala 29:58]
  assign _T_1015 = _T_1007[1:0]; // @[LZD.scala 44:32]
  assign _T_1016 = _T_1015 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1017 = _T_1015[1]; // @[LZD.scala 39:21]
  assign _T_1018 = _T_1015[0]; // @[LZD.scala 39:30]
  assign _T_1019 = ~ _T_1018; // @[LZD.scala 39:27]
  assign _T_1020 = _T_1017 | _T_1019; // @[LZD.scala 39:25]
  assign _T_1021 = {_T_1016,_T_1020}; // @[Cat.scala 29:58]
  assign _T_1022 = _T_1014[1]; // @[Shift.scala 12:21]
  assign _T_1023 = _T_1021[1]; // @[Shift.scala 12:21]
  assign _T_1024 = _T_1022 | _T_1023; // @[LZD.scala 49:16]
  assign _T_1025 = ~ _T_1023; // @[LZD.scala 49:27]
  assign _T_1026 = _T_1022 | _T_1025; // @[LZD.scala 49:25]
  assign _T_1027 = _T_1014[0:0]; // @[LZD.scala 49:47]
  assign _T_1028 = _T_1021[0:0]; // @[LZD.scala 49:59]
  assign _T_1029 = _T_1022 ? _T_1027 : _T_1028; // @[LZD.scala 49:35]
  assign _T_1031 = {_T_1024,_T_1026,_T_1029}; // @[Cat.scala 29:58]
  assign _T_1032 = _T_1006[2]; // @[Shift.scala 12:21]
  assign _T_1033 = _T_1031[2]; // @[Shift.scala 12:21]
  assign _T_1034 = _T_1032 | _T_1033; // @[LZD.scala 49:16]
  assign _T_1035 = ~ _T_1033; // @[LZD.scala 49:27]
  assign _T_1036 = _T_1032 | _T_1035; // @[LZD.scala 49:25]
  assign _T_1037 = _T_1006[1:0]; // @[LZD.scala 49:47]
  assign _T_1038 = _T_1031[1:0]; // @[LZD.scala 49:59]
  assign _T_1039 = _T_1032 ? _T_1037 : _T_1038; // @[LZD.scala 49:35]
  assign _T_1041 = {_T_1034,_T_1036,_T_1039}; // @[Cat.scala 29:58]
  assign _T_1042 = _T_980[7:0]; // @[LZD.scala 44:32]
  assign _T_1043 = _T_1042[7:4]; // @[LZD.scala 43:32]
  assign _T_1044 = _T_1043[3:2]; // @[LZD.scala 43:32]
  assign _T_1045 = _T_1044 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1046 = _T_1044[1]; // @[LZD.scala 39:21]
  assign _T_1047 = _T_1044[0]; // @[LZD.scala 39:30]
  assign _T_1048 = ~ _T_1047; // @[LZD.scala 39:27]
  assign _T_1049 = _T_1046 | _T_1048; // @[LZD.scala 39:25]
  assign _T_1050 = {_T_1045,_T_1049}; // @[Cat.scala 29:58]
  assign _T_1051 = _T_1043[1:0]; // @[LZD.scala 44:32]
  assign _T_1052 = _T_1051 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1053 = _T_1051[1]; // @[LZD.scala 39:21]
  assign _T_1054 = _T_1051[0]; // @[LZD.scala 39:30]
  assign _T_1055 = ~ _T_1054; // @[LZD.scala 39:27]
  assign _T_1056 = _T_1053 | _T_1055; // @[LZD.scala 39:25]
  assign _T_1057 = {_T_1052,_T_1056}; // @[Cat.scala 29:58]
  assign _T_1058 = _T_1050[1]; // @[Shift.scala 12:21]
  assign _T_1059 = _T_1057[1]; // @[Shift.scala 12:21]
  assign _T_1060 = _T_1058 | _T_1059; // @[LZD.scala 49:16]
  assign _T_1061 = ~ _T_1059; // @[LZD.scala 49:27]
  assign _T_1062 = _T_1058 | _T_1061; // @[LZD.scala 49:25]
  assign _T_1063 = _T_1050[0:0]; // @[LZD.scala 49:47]
  assign _T_1064 = _T_1057[0:0]; // @[LZD.scala 49:59]
  assign _T_1065 = _T_1058 ? _T_1063 : _T_1064; // @[LZD.scala 49:35]
  assign _T_1067 = {_T_1060,_T_1062,_T_1065}; // @[Cat.scala 29:58]
  assign _T_1068 = _T_1042[3:0]; // @[LZD.scala 44:32]
  assign _T_1069 = _T_1068[3:2]; // @[LZD.scala 43:32]
  assign _T_1070 = _T_1069 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1071 = _T_1069[1]; // @[LZD.scala 39:21]
  assign _T_1072 = _T_1069[0]; // @[LZD.scala 39:30]
  assign _T_1073 = ~ _T_1072; // @[LZD.scala 39:27]
  assign _T_1074 = _T_1071 | _T_1073; // @[LZD.scala 39:25]
  assign _T_1075 = {_T_1070,_T_1074}; // @[Cat.scala 29:58]
  assign _T_1076 = _T_1068[1:0]; // @[LZD.scala 44:32]
  assign _T_1077 = _T_1076 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1078 = _T_1076[1]; // @[LZD.scala 39:21]
  assign _T_1079 = _T_1076[0]; // @[LZD.scala 39:30]
  assign _T_1080 = ~ _T_1079; // @[LZD.scala 39:27]
  assign _T_1081 = _T_1078 | _T_1080; // @[LZD.scala 39:25]
  assign _T_1082 = {_T_1077,_T_1081}; // @[Cat.scala 29:58]
  assign _T_1083 = _T_1075[1]; // @[Shift.scala 12:21]
  assign _T_1084 = _T_1082[1]; // @[Shift.scala 12:21]
  assign _T_1085 = _T_1083 | _T_1084; // @[LZD.scala 49:16]
  assign _T_1086 = ~ _T_1084; // @[LZD.scala 49:27]
  assign _T_1087 = _T_1083 | _T_1086; // @[LZD.scala 49:25]
  assign _T_1088 = _T_1075[0:0]; // @[LZD.scala 49:47]
  assign _T_1089 = _T_1082[0:0]; // @[LZD.scala 49:59]
  assign _T_1090 = _T_1083 ? _T_1088 : _T_1089; // @[LZD.scala 49:35]
  assign _T_1092 = {_T_1085,_T_1087,_T_1090}; // @[Cat.scala 29:58]
  assign _T_1093 = _T_1067[2]; // @[Shift.scala 12:21]
  assign _T_1094 = _T_1092[2]; // @[Shift.scala 12:21]
  assign _T_1095 = _T_1093 | _T_1094; // @[LZD.scala 49:16]
  assign _T_1096 = ~ _T_1094; // @[LZD.scala 49:27]
  assign _T_1097 = _T_1093 | _T_1096; // @[LZD.scala 49:25]
  assign _T_1098 = _T_1067[1:0]; // @[LZD.scala 49:47]
  assign _T_1099 = _T_1092[1:0]; // @[LZD.scala 49:59]
  assign _T_1100 = _T_1093 ? _T_1098 : _T_1099; // @[LZD.scala 49:35]
  assign _T_1102 = {_T_1095,_T_1097,_T_1100}; // @[Cat.scala 29:58]
  assign _T_1103 = _T_1041[3]; // @[Shift.scala 12:21]
  assign _T_1104 = _T_1102[3]; // @[Shift.scala 12:21]
  assign _T_1105 = _T_1103 | _T_1104; // @[LZD.scala 49:16]
  assign _T_1106 = ~ _T_1104; // @[LZD.scala 49:27]
  assign _T_1107 = _T_1103 | _T_1106; // @[LZD.scala 49:25]
  assign _T_1108 = _T_1041[2:0]; // @[LZD.scala 49:47]
  assign _T_1109 = _T_1102[2:0]; // @[LZD.scala 49:59]
  assign _T_1110 = _T_1103 ? _T_1108 : _T_1109; // @[LZD.scala 49:35]
  assign _T_1112 = {_T_1105,_T_1107,_T_1110}; // @[Cat.scala 29:58]
  assign _T_1113 = _T_979[15:0]; // @[LZD.scala 44:32]
  assign _T_1114 = _T_1113[15:8]; // @[LZD.scala 43:32]
  assign _T_1115 = _T_1114[7:4]; // @[LZD.scala 43:32]
  assign _T_1116 = _T_1115[3:2]; // @[LZD.scala 43:32]
  assign _T_1117 = _T_1116 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1118 = _T_1116[1]; // @[LZD.scala 39:21]
  assign _T_1119 = _T_1116[0]; // @[LZD.scala 39:30]
  assign _T_1120 = ~ _T_1119; // @[LZD.scala 39:27]
  assign _T_1121 = _T_1118 | _T_1120; // @[LZD.scala 39:25]
  assign _T_1122 = {_T_1117,_T_1121}; // @[Cat.scala 29:58]
  assign _T_1123 = _T_1115[1:0]; // @[LZD.scala 44:32]
  assign _T_1124 = _T_1123 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1125 = _T_1123[1]; // @[LZD.scala 39:21]
  assign _T_1126 = _T_1123[0]; // @[LZD.scala 39:30]
  assign _T_1127 = ~ _T_1126; // @[LZD.scala 39:27]
  assign _T_1128 = _T_1125 | _T_1127; // @[LZD.scala 39:25]
  assign _T_1129 = {_T_1124,_T_1128}; // @[Cat.scala 29:58]
  assign _T_1130 = _T_1122[1]; // @[Shift.scala 12:21]
  assign _T_1131 = _T_1129[1]; // @[Shift.scala 12:21]
  assign _T_1132 = _T_1130 | _T_1131; // @[LZD.scala 49:16]
  assign _T_1133 = ~ _T_1131; // @[LZD.scala 49:27]
  assign _T_1134 = _T_1130 | _T_1133; // @[LZD.scala 49:25]
  assign _T_1135 = _T_1122[0:0]; // @[LZD.scala 49:47]
  assign _T_1136 = _T_1129[0:0]; // @[LZD.scala 49:59]
  assign _T_1137 = _T_1130 ? _T_1135 : _T_1136; // @[LZD.scala 49:35]
  assign _T_1139 = {_T_1132,_T_1134,_T_1137}; // @[Cat.scala 29:58]
  assign _T_1140 = _T_1114[3:0]; // @[LZD.scala 44:32]
  assign _T_1141 = _T_1140[3:2]; // @[LZD.scala 43:32]
  assign _T_1142 = _T_1141 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1143 = _T_1141[1]; // @[LZD.scala 39:21]
  assign _T_1144 = _T_1141[0]; // @[LZD.scala 39:30]
  assign _T_1145 = ~ _T_1144; // @[LZD.scala 39:27]
  assign _T_1146 = _T_1143 | _T_1145; // @[LZD.scala 39:25]
  assign _T_1147 = {_T_1142,_T_1146}; // @[Cat.scala 29:58]
  assign _T_1148 = _T_1140[1:0]; // @[LZD.scala 44:32]
  assign _T_1149 = _T_1148 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1150 = _T_1148[1]; // @[LZD.scala 39:21]
  assign _T_1151 = _T_1148[0]; // @[LZD.scala 39:30]
  assign _T_1152 = ~ _T_1151; // @[LZD.scala 39:27]
  assign _T_1153 = _T_1150 | _T_1152; // @[LZD.scala 39:25]
  assign _T_1154 = {_T_1149,_T_1153}; // @[Cat.scala 29:58]
  assign _T_1155 = _T_1147[1]; // @[Shift.scala 12:21]
  assign _T_1156 = _T_1154[1]; // @[Shift.scala 12:21]
  assign _T_1157 = _T_1155 | _T_1156; // @[LZD.scala 49:16]
  assign _T_1158 = ~ _T_1156; // @[LZD.scala 49:27]
  assign _T_1159 = _T_1155 | _T_1158; // @[LZD.scala 49:25]
  assign _T_1160 = _T_1147[0:0]; // @[LZD.scala 49:47]
  assign _T_1161 = _T_1154[0:0]; // @[LZD.scala 49:59]
  assign _T_1162 = _T_1155 ? _T_1160 : _T_1161; // @[LZD.scala 49:35]
  assign _T_1164 = {_T_1157,_T_1159,_T_1162}; // @[Cat.scala 29:58]
  assign _T_1165 = _T_1139[2]; // @[Shift.scala 12:21]
  assign _T_1166 = _T_1164[2]; // @[Shift.scala 12:21]
  assign _T_1167 = _T_1165 | _T_1166; // @[LZD.scala 49:16]
  assign _T_1168 = ~ _T_1166; // @[LZD.scala 49:27]
  assign _T_1169 = _T_1165 | _T_1168; // @[LZD.scala 49:25]
  assign _T_1170 = _T_1139[1:0]; // @[LZD.scala 49:47]
  assign _T_1171 = _T_1164[1:0]; // @[LZD.scala 49:59]
  assign _T_1172 = _T_1165 ? _T_1170 : _T_1171; // @[LZD.scala 49:35]
  assign _T_1174 = {_T_1167,_T_1169,_T_1172}; // @[Cat.scala 29:58]
  assign _T_1175 = _T_1113[7:0]; // @[LZD.scala 44:32]
  assign _T_1176 = _T_1175[7:4]; // @[LZD.scala 43:32]
  assign _T_1177 = _T_1176[3:2]; // @[LZD.scala 43:32]
  assign _T_1178 = _T_1177 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1179 = _T_1177[1]; // @[LZD.scala 39:21]
  assign _T_1180 = _T_1177[0]; // @[LZD.scala 39:30]
  assign _T_1181 = ~ _T_1180; // @[LZD.scala 39:27]
  assign _T_1182 = _T_1179 | _T_1181; // @[LZD.scala 39:25]
  assign _T_1183 = {_T_1178,_T_1182}; // @[Cat.scala 29:58]
  assign _T_1184 = _T_1176[1:0]; // @[LZD.scala 44:32]
  assign _T_1185 = _T_1184 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1186 = _T_1184[1]; // @[LZD.scala 39:21]
  assign _T_1187 = _T_1184[0]; // @[LZD.scala 39:30]
  assign _T_1188 = ~ _T_1187; // @[LZD.scala 39:27]
  assign _T_1189 = _T_1186 | _T_1188; // @[LZD.scala 39:25]
  assign _T_1190 = {_T_1185,_T_1189}; // @[Cat.scala 29:58]
  assign _T_1191 = _T_1183[1]; // @[Shift.scala 12:21]
  assign _T_1192 = _T_1190[1]; // @[Shift.scala 12:21]
  assign _T_1193 = _T_1191 | _T_1192; // @[LZD.scala 49:16]
  assign _T_1194 = ~ _T_1192; // @[LZD.scala 49:27]
  assign _T_1195 = _T_1191 | _T_1194; // @[LZD.scala 49:25]
  assign _T_1196 = _T_1183[0:0]; // @[LZD.scala 49:47]
  assign _T_1197 = _T_1190[0:0]; // @[LZD.scala 49:59]
  assign _T_1198 = _T_1191 ? _T_1196 : _T_1197; // @[LZD.scala 49:35]
  assign _T_1200 = {_T_1193,_T_1195,_T_1198}; // @[Cat.scala 29:58]
  assign _T_1201 = _T_1175[3:0]; // @[LZD.scala 44:32]
  assign _T_1202 = _T_1201[3:2]; // @[LZD.scala 43:32]
  assign _T_1203 = _T_1202 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1204 = _T_1202[1]; // @[LZD.scala 39:21]
  assign _T_1205 = _T_1202[0]; // @[LZD.scala 39:30]
  assign _T_1206 = ~ _T_1205; // @[LZD.scala 39:27]
  assign _T_1207 = _T_1204 | _T_1206; // @[LZD.scala 39:25]
  assign _T_1208 = {_T_1203,_T_1207}; // @[Cat.scala 29:58]
  assign _T_1209 = _T_1201[1:0]; // @[LZD.scala 44:32]
  assign _T_1210 = _T_1209 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1211 = _T_1209[1]; // @[LZD.scala 39:21]
  assign _T_1212 = _T_1209[0]; // @[LZD.scala 39:30]
  assign _T_1213 = ~ _T_1212; // @[LZD.scala 39:27]
  assign _T_1214 = _T_1211 | _T_1213; // @[LZD.scala 39:25]
  assign _T_1215 = {_T_1210,_T_1214}; // @[Cat.scala 29:58]
  assign _T_1216 = _T_1208[1]; // @[Shift.scala 12:21]
  assign _T_1217 = _T_1215[1]; // @[Shift.scala 12:21]
  assign _T_1218 = _T_1216 | _T_1217; // @[LZD.scala 49:16]
  assign _T_1219 = ~ _T_1217; // @[LZD.scala 49:27]
  assign _T_1220 = _T_1216 | _T_1219; // @[LZD.scala 49:25]
  assign _T_1221 = _T_1208[0:0]; // @[LZD.scala 49:47]
  assign _T_1222 = _T_1215[0:0]; // @[LZD.scala 49:59]
  assign _T_1223 = _T_1216 ? _T_1221 : _T_1222; // @[LZD.scala 49:35]
  assign _T_1225 = {_T_1218,_T_1220,_T_1223}; // @[Cat.scala 29:58]
  assign _T_1226 = _T_1200[2]; // @[Shift.scala 12:21]
  assign _T_1227 = _T_1225[2]; // @[Shift.scala 12:21]
  assign _T_1228 = _T_1226 | _T_1227; // @[LZD.scala 49:16]
  assign _T_1229 = ~ _T_1227; // @[LZD.scala 49:27]
  assign _T_1230 = _T_1226 | _T_1229; // @[LZD.scala 49:25]
  assign _T_1231 = _T_1200[1:0]; // @[LZD.scala 49:47]
  assign _T_1232 = _T_1225[1:0]; // @[LZD.scala 49:59]
  assign _T_1233 = _T_1226 ? _T_1231 : _T_1232; // @[LZD.scala 49:35]
  assign _T_1235 = {_T_1228,_T_1230,_T_1233}; // @[Cat.scala 29:58]
  assign _T_1236 = _T_1174[3]; // @[Shift.scala 12:21]
  assign _T_1237 = _T_1235[3]; // @[Shift.scala 12:21]
  assign _T_1238 = _T_1236 | _T_1237; // @[LZD.scala 49:16]
  assign _T_1239 = ~ _T_1237; // @[LZD.scala 49:27]
  assign _T_1240 = _T_1236 | _T_1239; // @[LZD.scala 49:25]
  assign _T_1241 = _T_1174[2:0]; // @[LZD.scala 49:47]
  assign _T_1242 = _T_1235[2:0]; // @[LZD.scala 49:59]
  assign _T_1243 = _T_1236 ? _T_1241 : _T_1242; // @[LZD.scala 49:35]
  assign _T_1245 = {_T_1238,_T_1240,_T_1243}; // @[Cat.scala 29:58]
  assign _T_1246 = _T_1112[4]; // @[Shift.scala 12:21]
  assign _T_1247 = _T_1245[4]; // @[Shift.scala 12:21]
  assign _T_1248 = _T_1246 | _T_1247; // @[LZD.scala 49:16]
  assign _T_1249 = ~ _T_1247; // @[LZD.scala 49:27]
  assign _T_1250 = _T_1246 | _T_1249; // @[LZD.scala 49:25]
  assign _T_1251 = _T_1112[3:0]; // @[LZD.scala 49:47]
  assign _T_1252 = _T_1245[3:0]; // @[LZD.scala 49:59]
  assign _T_1253 = _T_1246 ? _T_1251 : _T_1252; // @[LZD.scala 49:35]
  assign _T_1255 = {_T_1248,_T_1250,_T_1253}; // @[Cat.scala 29:58]
  assign _T_1256 = sumXor[14:0]; // @[LZD.scala 44:32]
  assign _T_1257 = _T_1256[14:7]; // @[LZD.scala 43:32]
  assign _T_1258 = _T_1257[7:4]; // @[LZD.scala 43:32]
  assign _T_1259 = _T_1258[3:2]; // @[LZD.scala 43:32]
  assign _T_1260 = _T_1259 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1261 = _T_1259[1]; // @[LZD.scala 39:21]
  assign _T_1262 = _T_1259[0]; // @[LZD.scala 39:30]
  assign _T_1263 = ~ _T_1262; // @[LZD.scala 39:27]
  assign _T_1264 = _T_1261 | _T_1263; // @[LZD.scala 39:25]
  assign _T_1265 = {_T_1260,_T_1264}; // @[Cat.scala 29:58]
  assign _T_1266 = _T_1258[1:0]; // @[LZD.scala 44:32]
  assign _T_1267 = _T_1266 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1268 = _T_1266[1]; // @[LZD.scala 39:21]
  assign _T_1269 = _T_1266[0]; // @[LZD.scala 39:30]
  assign _T_1270 = ~ _T_1269; // @[LZD.scala 39:27]
  assign _T_1271 = _T_1268 | _T_1270; // @[LZD.scala 39:25]
  assign _T_1272 = {_T_1267,_T_1271}; // @[Cat.scala 29:58]
  assign _T_1273 = _T_1265[1]; // @[Shift.scala 12:21]
  assign _T_1274 = _T_1272[1]; // @[Shift.scala 12:21]
  assign _T_1275 = _T_1273 | _T_1274; // @[LZD.scala 49:16]
  assign _T_1276 = ~ _T_1274; // @[LZD.scala 49:27]
  assign _T_1277 = _T_1273 | _T_1276; // @[LZD.scala 49:25]
  assign _T_1278 = _T_1265[0:0]; // @[LZD.scala 49:47]
  assign _T_1279 = _T_1272[0:0]; // @[LZD.scala 49:59]
  assign _T_1280 = _T_1273 ? _T_1278 : _T_1279; // @[LZD.scala 49:35]
  assign _T_1282 = {_T_1275,_T_1277,_T_1280}; // @[Cat.scala 29:58]
  assign _T_1283 = _T_1257[3:0]; // @[LZD.scala 44:32]
  assign _T_1284 = _T_1283[3:2]; // @[LZD.scala 43:32]
  assign _T_1285 = _T_1284 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1286 = _T_1284[1]; // @[LZD.scala 39:21]
  assign _T_1287 = _T_1284[0]; // @[LZD.scala 39:30]
  assign _T_1288 = ~ _T_1287; // @[LZD.scala 39:27]
  assign _T_1289 = _T_1286 | _T_1288; // @[LZD.scala 39:25]
  assign _T_1290 = {_T_1285,_T_1289}; // @[Cat.scala 29:58]
  assign _T_1291 = _T_1283[1:0]; // @[LZD.scala 44:32]
  assign _T_1292 = _T_1291 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1293 = _T_1291[1]; // @[LZD.scala 39:21]
  assign _T_1294 = _T_1291[0]; // @[LZD.scala 39:30]
  assign _T_1295 = ~ _T_1294; // @[LZD.scala 39:27]
  assign _T_1296 = _T_1293 | _T_1295; // @[LZD.scala 39:25]
  assign _T_1297 = {_T_1292,_T_1296}; // @[Cat.scala 29:58]
  assign _T_1298 = _T_1290[1]; // @[Shift.scala 12:21]
  assign _T_1299 = _T_1297[1]; // @[Shift.scala 12:21]
  assign _T_1300 = _T_1298 | _T_1299; // @[LZD.scala 49:16]
  assign _T_1301 = ~ _T_1299; // @[LZD.scala 49:27]
  assign _T_1302 = _T_1298 | _T_1301; // @[LZD.scala 49:25]
  assign _T_1303 = _T_1290[0:0]; // @[LZD.scala 49:47]
  assign _T_1304 = _T_1297[0:0]; // @[LZD.scala 49:59]
  assign _T_1305 = _T_1298 ? _T_1303 : _T_1304; // @[LZD.scala 49:35]
  assign _T_1307 = {_T_1300,_T_1302,_T_1305}; // @[Cat.scala 29:58]
  assign _T_1308 = _T_1282[2]; // @[Shift.scala 12:21]
  assign _T_1309 = _T_1307[2]; // @[Shift.scala 12:21]
  assign _T_1310 = _T_1308 | _T_1309; // @[LZD.scala 49:16]
  assign _T_1311 = ~ _T_1309; // @[LZD.scala 49:27]
  assign _T_1312 = _T_1308 | _T_1311; // @[LZD.scala 49:25]
  assign _T_1313 = _T_1282[1:0]; // @[LZD.scala 49:47]
  assign _T_1314 = _T_1307[1:0]; // @[LZD.scala 49:59]
  assign _T_1315 = _T_1308 ? _T_1313 : _T_1314; // @[LZD.scala 49:35]
  assign _T_1317 = {_T_1310,_T_1312,_T_1315}; // @[Cat.scala 29:58]
  assign _T_1318 = _T_1256[6:0]; // @[LZD.scala 44:32]
  assign _T_1319 = _T_1318[6:3]; // @[LZD.scala 43:32]
  assign _T_1320 = _T_1319[3:2]; // @[LZD.scala 43:32]
  assign _T_1321 = _T_1320 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1322 = _T_1320[1]; // @[LZD.scala 39:21]
  assign _T_1323 = _T_1320[0]; // @[LZD.scala 39:30]
  assign _T_1324 = ~ _T_1323; // @[LZD.scala 39:27]
  assign _T_1325 = _T_1322 | _T_1324; // @[LZD.scala 39:25]
  assign _T_1326 = {_T_1321,_T_1325}; // @[Cat.scala 29:58]
  assign _T_1327 = _T_1319[1:0]; // @[LZD.scala 44:32]
  assign _T_1328 = _T_1327 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1329 = _T_1327[1]; // @[LZD.scala 39:21]
  assign _T_1330 = _T_1327[0]; // @[LZD.scala 39:30]
  assign _T_1331 = ~ _T_1330; // @[LZD.scala 39:27]
  assign _T_1332 = _T_1329 | _T_1331; // @[LZD.scala 39:25]
  assign _T_1333 = {_T_1328,_T_1332}; // @[Cat.scala 29:58]
  assign _T_1334 = _T_1326[1]; // @[Shift.scala 12:21]
  assign _T_1335 = _T_1333[1]; // @[Shift.scala 12:21]
  assign _T_1336 = _T_1334 | _T_1335; // @[LZD.scala 49:16]
  assign _T_1337 = ~ _T_1335; // @[LZD.scala 49:27]
  assign _T_1338 = _T_1334 | _T_1337; // @[LZD.scala 49:25]
  assign _T_1339 = _T_1326[0:0]; // @[LZD.scala 49:47]
  assign _T_1340 = _T_1333[0:0]; // @[LZD.scala 49:59]
  assign _T_1341 = _T_1334 ? _T_1339 : _T_1340; // @[LZD.scala 49:35]
  assign _T_1343 = {_T_1336,_T_1338,_T_1341}; // @[Cat.scala 29:58]
  assign _T_1344 = _T_1318[2:0]; // @[LZD.scala 44:32]
  assign _T_1345 = _T_1344[2:1]; // @[LZD.scala 43:32]
  assign _T_1346 = _T_1345 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1347 = _T_1345[1]; // @[LZD.scala 39:21]
  assign _T_1348 = _T_1345[0]; // @[LZD.scala 39:30]
  assign _T_1349 = ~ _T_1348; // @[LZD.scala 39:27]
  assign _T_1350 = _T_1347 | _T_1349; // @[LZD.scala 39:25]
  assign _T_1351 = {_T_1346,_T_1350}; // @[Cat.scala 29:58]
  assign _T_1352 = _T_1344[0:0]; // @[LZD.scala 44:32]
  assign _T_1354 = _T_1351[1]; // @[Shift.scala 12:21]
  assign _T_1356 = _T_1351[0:0]; // @[LZD.scala 55:32]
  assign _T_1357 = _T_1354 ? _T_1356 : _T_1352; // @[LZD.scala 55:20]
  assign _T_1358 = {_T_1354,_T_1357}; // @[Cat.scala 29:58]
  assign _T_1359 = _T_1343[2]; // @[Shift.scala 12:21]
  assign _T_1361 = _T_1343[1:0]; // @[LZD.scala 55:32]
  assign _T_1362 = _T_1359 ? _T_1361 : _T_1358; // @[LZD.scala 55:20]
  assign _T_1363 = {_T_1359,_T_1362}; // @[Cat.scala 29:58]
  assign _T_1364 = _T_1317[3]; // @[Shift.scala 12:21]
  assign _T_1366 = _T_1317[2:0]; // @[LZD.scala 55:32]
  assign _T_1367 = _T_1364 ? _T_1366 : _T_1363; // @[LZD.scala 55:20]
  assign _T_1369 = _T_1255[5]; // @[Shift.scala 12:21]
  assign _T_1371 = {1'h1,_T_1364,_T_1367}; // @[Cat.scala 29:58]
  assign _T_1372 = _T_1255[4:0]; // @[LZD.scala 55:32]
  assign _T_1373 = _T_1369 ? _T_1372 : _T_1371; // @[LZD.scala 55:20]
  assign sumLZD = {_T_1369,_T_1373}; // @[Cat.scala 29:58]
  assign shiftValue = ~ sumLZD; // @[PositFMA.scala 126:24]
  assign _T_1374 = signSumSig[45:0]; // @[PositFMA.scala 127:38]
  assign _T_1375 = shiftValue < 6'h2e; // @[Shift.scala 16:24]
  assign _T_1377 = shiftValue[5]; // @[Shift.scala 12:21]
  assign _T_1378 = _T_1374[13:0]; // @[Shift.scala 64:52]
  assign _T_1380 = {_T_1378,32'h0}; // @[Cat.scala 29:58]
  assign _T_1381 = _T_1377 ? _T_1380 : _T_1374; // @[Shift.scala 64:27]
  assign _T_1382 = shiftValue[4:0]; // @[Shift.scala 66:70]
  assign _T_1383 = _T_1382[4]; // @[Shift.scala 12:21]
  assign _T_1384 = _T_1381[29:0]; // @[Shift.scala 64:52]
  assign _T_1386 = {_T_1384,16'h0}; // @[Cat.scala 29:58]
  assign _T_1387 = _T_1383 ? _T_1386 : _T_1381; // @[Shift.scala 64:27]
  assign _T_1388 = _T_1382[3:0]; // @[Shift.scala 66:70]
  assign _T_1389 = _T_1388[3]; // @[Shift.scala 12:21]
  assign _T_1390 = _T_1387[37:0]; // @[Shift.scala 64:52]
  assign _T_1392 = {_T_1390,8'h0}; // @[Cat.scala 29:58]
  assign _T_1393 = _T_1389 ? _T_1392 : _T_1387; // @[Shift.scala 64:27]
  assign _T_1394 = _T_1388[2:0]; // @[Shift.scala 66:70]
  assign _T_1395 = _T_1394[2]; // @[Shift.scala 12:21]
  assign _T_1396 = _T_1393[41:0]; // @[Shift.scala 64:52]
  assign _T_1398 = {_T_1396,4'h0}; // @[Cat.scala 29:58]
  assign _T_1399 = _T_1395 ? _T_1398 : _T_1393; // @[Shift.scala 64:27]
  assign _T_1400 = _T_1394[1:0]; // @[Shift.scala 66:70]
  assign _T_1401 = _T_1400[1]; // @[Shift.scala 12:21]
  assign _T_1402 = _T_1399[43:0]; // @[Shift.scala 64:52]
  assign _T_1404 = {_T_1402,2'h0}; // @[Cat.scala 29:58]
  assign _T_1405 = _T_1401 ? _T_1404 : _T_1399; // @[Shift.scala 64:27]
  assign _T_1406 = _T_1400[0:0]; // @[Shift.scala 66:70]
  assign _T_1408 = _T_1405[44:0]; // @[Shift.scala 64:52]
  assign _T_1409 = {_T_1408,1'h0}; // @[Cat.scala 29:58]
  assign _T_1410 = _T_1406 ? _T_1409 : _T_1405; // @[Shift.scala 64:27]
  assign normalFracTmp = _T_1375 ? _T_1410 : 46'h0; // @[Shift.scala 16:10]
  assign _T_1412 = $signed(greaterScale) + $signed(10'sh2); // @[PositFMA.scala 130:36]
  assign _T_1413 = $signed(_T_1412); // @[PositFMA.scala 130:36]
  assign _T_1414 = {1'h1,_T_1369,_T_1373}; // @[Cat.scala 29:58]
  assign _T_1415 = $signed(_T_1414); // @[PositFMA.scala 130:61]
  assign _GEN_20 = {{3{_T_1415[6]}},_T_1415}; // @[PositFMA.scala 130:42]
  assign _T_1417 = $signed(_T_1413) + $signed(_GEN_20); // @[PositFMA.scala 130:42]
  assign sumScale = $signed(_T_1417); // @[PositFMA.scala 130:42]
  assign sumFrac = normalFracTmp[45:24]; // @[PositFMA.scala 131:41]
  assign grsTmp = normalFracTmp[23:0]; // @[PositFMA.scala 134:41]
  assign _T_1418 = grsTmp[23:22]; // @[PositFMA.scala 137:40]
  assign _T_1419 = grsTmp[21:0]; // @[PositFMA.scala 137:56]
  assign _T_1420 = _T_1419 != 22'h0; // @[PositFMA.scala 137:60]
  assign underflow = $signed(sumScale) < $signed(-10'shd1); // @[PositFMA.scala 144:32]
  assign overflow = $signed(sumScale) > $signed(10'shd0); // @[PositFMA.scala 145:32]
  assign _T_1421 = signSumSig != 48'h0; // @[PositFMA.scala 154:32]
  assign decF_isZero = ~ _T_1421; // @[PositFMA.scala 154:20]
  assign _T_1423 = underflow ? $signed(-10'shd1) : $signed(sumScale); // @[Mux.scala 87:16]
  assign _T_1424 = overflow ? $signed(10'shd0) : $signed(_T_1423); // @[Mux.scala 87:16]
  assign _GEN_21 = _T_1424[8:0]; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  assign decF_scale = $signed(_GEN_21); // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  assign _T_1425 = decF_scale[2:0]; // @[convert.scala 46:61]
  assign _T_1426 = ~ _T_1425; // @[convert.scala 46:52]
  assign _T_1428 = sumSign ? _T_1426 : _T_1425; // @[convert.scala 46:42]
  assign _T_1429 = decF_scale[8:3]; // @[convert.scala 48:34]
  assign _T_1430 = _T_1429[5:5]; // @[convert.scala 49:36]
  assign _T_1432 = ~ _T_1429; // @[convert.scala 50:36]
  assign _T_1433 = $signed(_T_1432); // @[convert.scala 50:36]
  assign _T_1434 = _T_1430 ? $signed(_T_1433) : $signed(_T_1429); // @[convert.scala 50:28]
  assign _T_1435 = _T_1430 ^ sumSign; // @[convert.scala 51:31]
  assign _T_1436 = ~ _T_1435; // @[convert.scala 52:43]
  assign _T_1440 = {_T_1436,_T_1435,_T_1428,sumFrac,_T_1418,_T_1420}; // @[Cat.scala 29:58]
  assign _T_1441 = $unsigned(_T_1434); // @[Shift.scala 39:17]
  assign _T_1442 = _T_1441 < 6'h1e; // @[Shift.scala 39:24]
  assign _T_1443 = _T_1434[4:0]; // @[Shift.scala 40:44]
  assign _T_1444 = _T_1440[29:16]; // @[Shift.scala 90:30]
  assign _T_1445 = _T_1440[15:0]; // @[Shift.scala 90:48]
  assign _T_1446 = _T_1445 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_22 = {{13'd0}, _T_1446}; // @[Shift.scala 90:39]
  assign _T_1447 = _T_1444 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_1448 = _T_1443[4]; // @[Shift.scala 12:21]
  assign _T_1449 = _T_1440[29]; // @[Shift.scala 12:21]
  assign _T_1451 = _T_1449 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_1452 = {_T_1451,_T_1447}; // @[Cat.scala 29:58]
  assign _T_1453 = _T_1448 ? _T_1452 : _T_1440; // @[Shift.scala 91:22]
  assign _T_1454 = _T_1443[3:0]; // @[Shift.scala 92:77]
  assign _T_1455 = _T_1453[29:8]; // @[Shift.scala 90:30]
  assign _T_1456 = _T_1453[7:0]; // @[Shift.scala 90:48]
  assign _T_1457 = _T_1456 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_23 = {{21'd0}, _T_1457}; // @[Shift.scala 90:39]
  assign _T_1458 = _T_1455 | _GEN_23; // @[Shift.scala 90:39]
  assign _T_1459 = _T_1454[3]; // @[Shift.scala 12:21]
  assign _T_1460 = _T_1453[29]; // @[Shift.scala 12:21]
  assign _T_1462 = _T_1460 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_1463 = {_T_1462,_T_1458}; // @[Cat.scala 29:58]
  assign _T_1464 = _T_1459 ? _T_1463 : _T_1453; // @[Shift.scala 91:22]
  assign _T_1465 = _T_1454[2:0]; // @[Shift.scala 92:77]
  assign _T_1466 = _T_1464[29:4]; // @[Shift.scala 90:30]
  assign _T_1467 = _T_1464[3:0]; // @[Shift.scala 90:48]
  assign _T_1468 = _T_1467 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_24 = {{25'd0}, _T_1468}; // @[Shift.scala 90:39]
  assign _T_1469 = _T_1466 | _GEN_24; // @[Shift.scala 90:39]
  assign _T_1470 = _T_1465[2]; // @[Shift.scala 12:21]
  assign _T_1471 = _T_1464[29]; // @[Shift.scala 12:21]
  assign _T_1473 = _T_1471 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_1474 = {_T_1473,_T_1469}; // @[Cat.scala 29:58]
  assign _T_1475 = _T_1470 ? _T_1474 : _T_1464; // @[Shift.scala 91:22]
  assign _T_1476 = _T_1465[1:0]; // @[Shift.scala 92:77]
  assign _T_1477 = _T_1475[29:2]; // @[Shift.scala 90:30]
  assign _T_1478 = _T_1475[1:0]; // @[Shift.scala 90:48]
  assign _T_1479 = _T_1478 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_25 = {{27'd0}, _T_1479}; // @[Shift.scala 90:39]
  assign _T_1480 = _T_1477 | _GEN_25; // @[Shift.scala 90:39]
  assign _T_1481 = _T_1476[1]; // @[Shift.scala 12:21]
  assign _T_1482 = _T_1475[29]; // @[Shift.scala 12:21]
  assign _T_1484 = _T_1482 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_1485 = {_T_1484,_T_1480}; // @[Cat.scala 29:58]
  assign _T_1486 = _T_1481 ? _T_1485 : _T_1475; // @[Shift.scala 91:22]
  assign _T_1487 = _T_1476[0:0]; // @[Shift.scala 92:77]
  assign _T_1488 = _T_1486[29:1]; // @[Shift.scala 90:30]
  assign _T_1489 = _T_1486[0:0]; // @[Shift.scala 90:48]
  assign _GEN_26 = {{28'd0}, _T_1489}; // @[Shift.scala 90:39]
  assign _T_1491 = _T_1488 | _GEN_26; // @[Shift.scala 90:39]
  assign _T_1493 = _T_1486[29]; // @[Shift.scala 12:21]
  assign _T_1494 = {_T_1493,_T_1491}; // @[Cat.scala 29:58]
  assign _T_1495 = _T_1487 ? _T_1494 : _T_1486; // @[Shift.scala 91:22]
  assign _T_1498 = _T_1449 ? 30'h3fffffff : 30'h0; // @[Bitwise.scala 71:12]
  assign _T_1499 = _T_1442 ? _T_1495 : _T_1498; // @[Shift.scala 39:10]
  assign _T_1500 = _T_1499[3]; // @[convert.scala 55:31]
  assign _T_1501 = _T_1499[2]; // @[convert.scala 56:31]
  assign _T_1502 = _T_1499[1]; // @[convert.scala 57:31]
  assign _T_1503 = _T_1499[0]; // @[convert.scala 58:31]
  assign _T_1504 = _T_1499[29:3]; // @[convert.scala 59:69]
  assign _T_1505 = _T_1504 != 27'h0; // @[convert.scala 59:81]
  assign _T_1506 = ~ _T_1505; // @[convert.scala 59:50]
  assign _T_1508 = _T_1504 == 27'h7ffffff; // @[convert.scala 60:81]
  assign _T_1509 = _T_1500 | _T_1502; // @[convert.scala 61:44]
  assign _T_1510 = _T_1509 | _T_1503; // @[convert.scala 61:52]
  assign _T_1511 = _T_1501 & _T_1510; // @[convert.scala 61:36]
  assign _T_1512 = ~ _T_1508; // @[convert.scala 62:63]
  assign _T_1513 = _T_1512 & _T_1511; // @[convert.scala 62:103]
  assign _T_1514 = _T_1506 | _T_1513; // @[convert.scala 62:60]
  assign _GEN_27 = {{26'd0}, _T_1514}; // @[convert.scala 63:56]
  assign _T_1517 = _T_1504 + _GEN_27; // @[convert.scala 63:56]
  assign _T_1518 = {sumSign,_T_1517}; // @[Cat.scala 29:58]
  assign io_F = _T_1526; // @[PositFMA.scala 174:15]
  assign io_outValid = _T_1522; // @[PositFMA.scala 173:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  outIsNaR_phase2 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  mulSig_phase2 = _RAND_1[46:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  addFrac_phase2 = _RAND_2[21:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mulScale_phase2 = _RAND_3[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addScale_phase2 = _RAND_4[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addSign_phase2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addZero_phase2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  inValid_phase2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1522 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_1526 = _RAND_9[27:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (io_inValid) begin
      outIsNaR_phase2 <= outIsNaR;
    end
    if (io_inValid) begin
      mulSig_phase2 <= mulSig;
    end
    if (io_inValid) begin
      addFrac_phase2 <= decC_fraction;
    end
    if (io_inValid) begin
      mulScale_phase2 <= mulScale;
    end
    if (io_inValid) begin
      addScale_phase2 <= decC_scale;
    end
    if (io_inValid) begin
      addSign_phase2 <= _T_567;
    end
    if (io_inValid) begin
      addZero_phase2 <= decC_isZero;
    end
    if (reset) begin
      inValid_phase2 <= 1'h0;
    end else begin
      inValid_phase2 <= io_inValid;
    end
    if (reset) begin
      _T_1522 <= 1'h0;
    end else begin
      _T_1522 <= inValid_phase2;
    end
    if (inValid_phase2) begin
      if (outIsNaR_phase2) begin
        _T_1526 <= 28'h8000000;
      end else begin
        if (decF_isZero) begin
          _T_1526 <= 28'h0;
        end else begin
          _T_1526 <= _T_1518;
        end
      end
    end
  end
endmodule
