module PositDivSqrter12_1(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input  [11:0] io_A,
  input  [11:0] io_B,
  output        io_diviValid,
  output        io_sqrtValid,
  output        io_invalidExc,
  output [11:0] io_Q
);
  reg [3:0] cycleNum; // @[PositDivisionSqrt.scala 63:26]
  reg [31:0] _RAND_0;
  reg  sqrtOp_Z; // @[PositDivisionSqrt.scala 65:22]
  reg [31:0] _RAND_1;
  reg  isNaR_Z; // @[PositDivisionSqrt.scala 66:22]
  reg [31:0] _RAND_2;
  reg  isZero_Z; // @[PositDivisionSqrt.scala 67:22]
  reg [31:0] _RAND_3;
  reg [6:0] scale_Z; // @[PositDivisionSqrt.scala 68:22]
  reg [31:0] _RAND_4;
  reg  signB_Z; // @[PositDivisionSqrt.scala 69:28]
  reg [31:0] _RAND_5;
  reg [7:0] fractB_Z; // @[PositDivisionSqrt.scala 70:22]
  reg [31:0] _RAND_6;
  reg [14:0] rem_Z; // @[PositDivisionSqrt.scala 71:22]
  reg [31:0] _RAND_7;
  reg [14:0] sigX_Z; // @[PositDivisionSqrt.scala 72:22]
  reg [31:0] _RAND_8;
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [9:0] _T_4; // @[convert.scala 19:24]
  wire [9:0] _T_5; // @[convert.scala 19:43]
  wire [9:0] _T_6; // @[convert.scala 19:39]
  wire [7:0] _T_7; // @[LZD.scala 43:32]
  wire [3:0] _T_8; // @[LZD.scala 43:32]
  wire [1:0] _T_9; // @[LZD.scala 43:32]
  wire  _T_10; // @[LZD.scala 39:14]
  wire  _T_11; // @[LZD.scala 39:21]
  wire  _T_12; // @[LZD.scala 39:30]
  wire  _T_13; // @[LZD.scala 39:27]
  wire  _T_14; // @[LZD.scala 39:25]
  wire [1:0] _T_15; // @[Cat.scala 29:58]
  wire [1:0] _T_16; // @[LZD.scala 44:32]
  wire  _T_17; // @[LZD.scala 39:14]
  wire  _T_18; // @[LZD.scala 39:21]
  wire  _T_19; // @[LZD.scala 39:30]
  wire  _T_20; // @[LZD.scala 39:27]
  wire  _T_21; // @[LZD.scala 39:25]
  wire [1:0] _T_22; // @[Cat.scala 29:58]
  wire  _T_23; // @[Shift.scala 12:21]
  wire  _T_24; // @[Shift.scala 12:21]
  wire  _T_25; // @[LZD.scala 49:16]
  wire  _T_26; // @[LZD.scala 49:27]
  wire  _T_27; // @[LZD.scala 49:25]
  wire  _T_28; // @[LZD.scala 49:47]
  wire  _T_29; // @[LZD.scala 49:59]
  wire  _T_30; // @[LZD.scala 49:35]
  wire [2:0] _T_32; // @[Cat.scala 29:58]
  wire [3:0] _T_33; // @[LZD.scala 44:32]
  wire [1:0] _T_34; // @[LZD.scala 43:32]
  wire  _T_35; // @[LZD.scala 39:14]
  wire  _T_36; // @[LZD.scala 39:21]
  wire  _T_37; // @[LZD.scala 39:30]
  wire  _T_38; // @[LZD.scala 39:27]
  wire  _T_39; // @[LZD.scala 39:25]
  wire [1:0] _T_40; // @[Cat.scala 29:58]
  wire [1:0] _T_41; // @[LZD.scala 44:32]
  wire  _T_42; // @[LZD.scala 39:14]
  wire  _T_43; // @[LZD.scala 39:21]
  wire  _T_44; // @[LZD.scala 39:30]
  wire  _T_45; // @[LZD.scala 39:27]
  wire  _T_46; // @[LZD.scala 39:25]
  wire [1:0] _T_47; // @[Cat.scala 29:58]
  wire  _T_48; // @[Shift.scala 12:21]
  wire  _T_49; // @[Shift.scala 12:21]
  wire  _T_50; // @[LZD.scala 49:16]
  wire  _T_51; // @[LZD.scala 49:27]
  wire  _T_52; // @[LZD.scala 49:25]
  wire  _T_53; // @[LZD.scala 49:47]
  wire  _T_54; // @[LZD.scala 49:59]
  wire  _T_55; // @[LZD.scala 49:35]
  wire [2:0] _T_57; // @[Cat.scala 29:58]
  wire  _T_58; // @[Shift.scala 12:21]
  wire  _T_59; // @[Shift.scala 12:21]
  wire  _T_60; // @[LZD.scala 49:16]
  wire  _T_61; // @[LZD.scala 49:27]
  wire  _T_62; // @[LZD.scala 49:25]
  wire [1:0] _T_63; // @[LZD.scala 49:47]
  wire [1:0] _T_64; // @[LZD.scala 49:59]
  wire [1:0] _T_65; // @[LZD.scala 49:35]
  wire [3:0] _T_67; // @[Cat.scala 29:58]
  wire [1:0] _T_68; // @[LZD.scala 44:32]
  wire  _T_69; // @[LZD.scala 39:14]
  wire  _T_70; // @[LZD.scala 39:21]
  wire  _T_71; // @[LZD.scala 39:30]
  wire  _T_72; // @[LZD.scala 39:27]
  wire  _T_73; // @[LZD.scala 39:25]
  wire  _T_75; // @[Shift.scala 12:21]
  wire [2:0] _T_77; // @[Cat.scala 29:58]
  wire [2:0] _T_78; // @[LZD.scala 55:32]
  wire [2:0] _T_79; // @[LZD.scala 55:20]
  wire [3:0] _T_80; // @[Cat.scala 29:58]
  wire [3:0] _T_81; // @[convert.scala 21:22]
  wire [8:0] _T_82; // @[convert.scala 22:36]
  wire  _T_83; // @[Shift.scala 16:24]
  wire  _T_85; // @[Shift.scala 12:21]
  wire  _T_86; // @[Shift.scala 64:52]
  wire [8:0] _T_88; // @[Cat.scala 29:58]
  wire [8:0] _T_89; // @[Shift.scala 64:27]
  wire [2:0] _T_90; // @[Shift.scala 66:70]
  wire  _T_91; // @[Shift.scala 12:21]
  wire [4:0] _T_92; // @[Shift.scala 64:52]
  wire [8:0] _T_94; // @[Cat.scala 29:58]
  wire [8:0] _T_95; // @[Shift.scala 64:27]
  wire [1:0] _T_96; // @[Shift.scala 66:70]
  wire  _T_97; // @[Shift.scala 12:21]
  wire [6:0] _T_98; // @[Shift.scala 64:52]
  wire [8:0] _T_100; // @[Cat.scala 29:58]
  wire [8:0] _T_101; // @[Shift.scala 64:27]
  wire  _T_102; // @[Shift.scala 66:70]
  wire [7:0] _T_104; // @[Shift.scala 64:52]
  wire [8:0] _T_105; // @[Cat.scala 29:58]
  wire [8:0] _T_106; // @[Shift.scala 64:27]
  wire [8:0] _T_107; // @[Shift.scala 16:10]
  wire  _T_108; // @[convert.scala 23:34]
  wire [7:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_110; // @[convert.scala 25:26]
  wire [3:0] _T_112; // @[convert.scala 25:42]
  wire  _T_115; // @[convert.scala 26:67]
  wire  _T_116; // @[convert.scala 26:51]
  wire [5:0] _T_117; // @[Cat.scala 29:58]
  wire [10:0] _T_119; // @[convert.scala 29:56]
  wire  _T_120; // @[convert.scala 29:60]
  wire  _T_121; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_124; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [5:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_133; // @[convert.scala 18:24]
  wire  _T_134; // @[convert.scala 18:40]
  wire  _T_135; // @[convert.scala 18:36]
  wire [9:0] _T_136; // @[convert.scala 19:24]
  wire [9:0] _T_137; // @[convert.scala 19:43]
  wire [9:0] _T_138; // @[convert.scala 19:39]
  wire [7:0] _T_139; // @[LZD.scala 43:32]
  wire [3:0] _T_140; // @[LZD.scala 43:32]
  wire [1:0] _T_141; // @[LZD.scala 43:32]
  wire  _T_142; // @[LZD.scala 39:14]
  wire  _T_143; // @[LZD.scala 39:21]
  wire  _T_144; // @[LZD.scala 39:30]
  wire  _T_145; // @[LZD.scala 39:27]
  wire  _T_146; // @[LZD.scala 39:25]
  wire [1:0] _T_147; // @[Cat.scala 29:58]
  wire [1:0] _T_148; // @[LZD.scala 44:32]
  wire  _T_149; // @[LZD.scala 39:14]
  wire  _T_150; // @[LZD.scala 39:21]
  wire  _T_151; // @[LZD.scala 39:30]
  wire  _T_152; // @[LZD.scala 39:27]
  wire  _T_153; // @[LZD.scala 39:25]
  wire [1:0] _T_154; // @[Cat.scala 29:58]
  wire  _T_155; // @[Shift.scala 12:21]
  wire  _T_156; // @[Shift.scala 12:21]
  wire  _T_157; // @[LZD.scala 49:16]
  wire  _T_158; // @[LZD.scala 49:27]
  wire  _T_159; // @[LZD.scala 49:25]
  wire  _T_160; // @[LZD.scala 49:47]
  wire  _T_161; // @[LZD.scala 49:59]
  wire  _T_162; // @[LZD.scala 49:35]
  wire [2:0] _T_164; // @[Cat.scala 29:58]
  wire [3:0] _T_165; // @[LZD.scala 44:32]
  wire [1:0] _T_166; // @[LZD.scala 43:32]
  wire  _T_167; // @[LZD.scala 39:14]
  wire  _T_168; // @[LZD.scala 39:21]
  wire  _T_169; // @[LZD.scala 39:30]
  wire  _T_170; // @[LZD.scala 39:27]
  wire  _T_171; // @[LZD.scala 39:25]
  wire [1:0] _T_172; // @[Cat.scala 29:58]
  wire [1:0] _T_173; // @[LZD.scala 44:32]
  wire  _T_174; // @[LZD.scala 39:14]
  wire  _T_175; // @[LZD.scala 39:21]
  wire  _T_176; // @[LZD.scala 39:30]
  wire  _T_177; // @[LZD.scala 39:27]
  wire  _T_178; // @[LZD.scala 39:25]
  wire [1:0] _T_179; // @[Cat.scala 29:58]
  wire  _T_180; // @[Shift.scala 12:21]
  wire  _T_181; // @[Shift.scala 12:21]
  wire  _T_182; // @[LZD.scala 49:16]
  wire  _T_183; // @[LZD.scala 49:27]
  wire  _T_184; // @[LZD.scala 49:25]
  wire  _T_185; // @[LZD.scala 49:47]
  wire  _T_186; // @[LZD.scala 49:59]
  wire  _T_187; // @[LZD.scala 49:35]
  wire [2:0] _T_189; // @[Cat.scala 29:58]
  wire  _T_190; // @[Shift.scala 12:21]
  wire  _T_191; // @[Shift.scala 12:21]
  wire  _T_192; // @[LZD.scala 49:16]
  wire  _T_193; // @[LZD.scala 49:27]
  wire  _T_194; // @[LZD.scala 49:25]
  wire [1:0] _T_195; // @[LZD.scala 49:47]
  wire [1:0] _T_196; // @[LZD.scala 49:59]
  wire [1:0] _T_197; // @[LZD.scala 49:35]
  wire [3:0] _T_199; // @[Cat.scala 29:58]
  wire [1:0] _T_200; // @[LZD.scala 44:32]
  wire  _T_201; // @[LZD.scala 39:14]
  wire  _T_202; // @[LZD.scala 39:21]
  wire  _T_203; // @[LZD.scala 39:30]
  wire  _T_204; // @[LZD.scala 39:27]
  wire  _T_205; // @[LZD.scala 39:25]
  wire  _T_207; // @[Shift.scala 12:21]
  wire [2:0] _T_209; // @[Cat.scala 29:58]
  wire [2:0] _T_210; // @[LZD.scala 55:32]
  wire [2:0] _T_211; // @[LZD.scala 55:20]
  wire [3:0] _T_212; // @[Cat.scala 29:58]
  wire [3:0] _T_213; // @[convert.scala 21:22]
  wire [8:0] _T_214; // @[convert.scala 22:36]
  wire  _T_215; // @[Shift.scala 16:24]
  wire  _T_217; // @[Shift.scala 12:21]
  wire  _T_218; // @[Shift.scala 64:52]
  wire [8:0] _T_220; // @[Cat.scala 29:58]
  wire [8:0] _T_221; // @[Shift.scala 64:27]
  wire [2:0] _T_222; // @[Shift.scala 66:70]
  wire  _T_223; // @[Shift.scala 12:21]
  wire [4:0] _T_224; // @[Shift.scala 64:52]
  wire [8:0] _T_226; // @[Cat.scala 29:58]
  wire [8:0] _T_227; // @[Shift.scala 64:27]
  wire [1:0] _T_228; // @[Shift.scala 66:70]
  wire  _T_229; // @[Shift.scala 12:21]
  wire [6:0] _T_230; // @[Shift.scala 64:52]
  wire [8:0] _T_232; // @[Cat.scala 29:58]
  wire [8:0] _T_233; // @[Shift.scala 64:27]
  wire  _T_234; // @[Shift.scala 66:70]
  wire [7:0] _T_236; // @[Shift.scala 64:52]
  wire [8:0] _T_237; // @[Cat.scala 29:58]
  wire [8:0] _T_238; // @[Shift.scala 64:27]
  wire [8:0] _T_239; // @[Shift.scala 16:10]
  wire  _T_240; // @[convert.scala 23:34]
  wire [7:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_242; // @[convert.scala 25:26]
  wire [3:0] _T_244; // @[convert.scala 25:42]
  wire  _T_247; // @[convert.scala 26:67]
  wire  _T_248; // @[convert.scala 26:51]
  wire [5:0] _T_249; // @[Cat.scala 29:58]
  wire [10:0] _T_251; // @[convert.scala 29:56]
  wire  _T_252; // @[convert.scala 29:60]
  wire  _T_253; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_256; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [5:0] decB_scale; // @[convert.scala 32:24]
  wire [2:0] _T_265; // @[Bitwise.scala 71:12]
  wire  _T_266; // @[PositDivisionSqrt.scala 80:40]
  wire [14:0] sigA_S; // @[Cat.scala 29:58]
  wire  _T_269; // @[PositDivisionSqrt.scala 82:31]
  wire [14:0] sigB_S; // @[Cat.scala 29:58]
  wire  _T_272; // @[PositDivisionSqrt.scala 85:25]
  wire  invalidSqrt; // @[PositDivisionSqrt.scala 85:37]
  wire  _T_273; // @[PositDivisionSqrt.scala 88:42]
  wire  _T_274; // @[PositDivisionSqrt.scala 89:42]
  wire  _T_275; // @[PositDivisionSqrt.scala 89:56]
  wire  _T_276; // @[PositDivisionSqrt.scala 94:46]
  wire  _T_277; // @[PositDivisionSqrt.scala 94:43]
  wire  _T_278; // @[PositDivisionSqrt.scala 94:62]
  wire  _T_279; // @[PositDivisionSqrt.scala 94:59]
  wire  specialCaseA_S; // @[PositDivisionSqrt.scala 97:38]
  wire  specialCaseB_S; // @[PositDivisionSqrt.scala 98:38]
  wire  _T_280; // @[PositDivisionSqrt.scala 99:27]
  wire  _T_281; // @[PositDivisionSqrt.scala 99:46]
  wire  normalCase_S_div; // @[PositDivisionSqrt.scala 99:43]
  wire  normalCase_S_sqrt; // @[PositDivisionSqrt.scala 100:43]
  wire  normalCase_S; // @[PositDivisionSqrt.scala 101:30]
  wire [6:0] sExpQuot_S_div; // @[PositDivisionSqrt.scala 103:38]
  wire  _T_284; // @[PositDivisionSqrt.scala 104:50]
  wire  oddSqrt_S; // @[PositDivisionSqrt.scala 104:37]
  wire  idle; // @[PositDivisionSqrt.scala 109:39]
  wire  ready; // @[PositDivisionSqrt.scala 110:39]
  wire  entering; // @[PositDivisionSqrt.scala 111:35]
  wire  entering_normalCase; // @[PositDivisionSqrt.scala 112:38]
  wire  _T_285; // @[PositDivisionSqrt.scala 113:35]
  wire  _T_286; // @[PositDivisionSqrt.scala 113:58]
  wire  scaleNotChange; // @[PositDivisionSqrt.scala 113:50]
  wire  _T_287; // @[PositDivisionSqrt.scala 114:39]
  wire  skipCycle2; // @[PositDivisionSqrt.scala 114:48]
  wire  _T_288; // @[PositDivisionSqrt.scala 116:8]
  wire  _T_289; // @[PositDivisionSqrt.scala 116:14]
  wire  _T_290; // @[PositDivisionSqrt.scala 117:32]
  wire  _T_291; // @[PositDivisionSqrt.scala 117:30]
  wire [3:0] _T_293; // @[PositDivisionSqrt.scala 119:26]
  wire [3:0] _T_294; // @[PositDivisionSqrt.scala 118:20]
  wire [3:0] _GEN_9; // @[PositDivisionSqrt.scala 117:64]
  wire [3:0] _T_295; // @[PositDivisionSqrt.scala 117:64]
  wire  _T_297; // @[PositDivisionSqrt.scala 123:30]
  wire  _T_298; // @[PositDivisionSqrt.scala 123:27]
  wire [3:0] _T_300; // @[PositDivisionSqrt.scala 123:52]
  wire [3:0] _T_301; // @[PositDivisionSqrt.scala 123:20]
  wire [3:0] _T_302; // @[PositDivisionSqrt.scala 122:64]
  wire  _T_304; // @[PositDivisionSqrt.scala 124:27]
  wire [3:0] _GEN_10; // @[PositDivisionSqrt.scala 123:64]
  wire [3:0] _T_306; // @[PositDivisionSqrt.scala 123:64]
  wire [4:0] _T_307; // @[PositDivisionSqrt.scala 134:42]
  wire  _T_309; // @[PositDivisionSqrt.scala 137:31]
  wire  _T_310; // @[PositDivisionSqrt.scala 137:28]
  wire [15:0] _T_311; // @[PositDivisionSqrt.scala 146:22]
  wire [13:0] bitMask; // @[PositDivisionSqrt.scala 146:35]
  wire  _T_313; // @[PositDivisionSqrt.scala 148:26]
  wire  _T_314; // @[PositDivisionSqrt.scala 148:23]
  wire [14:0] _T_315; // @[PositDivisionSqrt.scala 148:16]
  wire  _T_316; // @[PositDivisionSqrt.scala 149:23]
  wire [15:0] _T_317; // @[PositDivisionSqrt.scala 149:46]
  wire [14:0] _T_318; // @[PositDivisionSqrt.scala 149:56]
  wire [14:0] _T_319; // @[PositDivisionSqrt.scala 149:16]
  wire [14:0] _T_320; // @[PositDivisionSqrt.scala 148:66]
  wire  _T_321; // @[PositDivisionSqrt.scala 150:17]
  wire [14:0] _T_322; // @[PositDivisionSqrt.scala 150:16]
  wire [14:0] rem; // @[PositDivisionSqrt.scala 149:66]
  wire  _T_324; // @[PositDivisionSqrt.scala 152:29]
  wire [14:0] _T_325; // @[PositDivisionSqrt.scala 152:22]
  wire  _T_326; // @[PositDivisionSqrt.scala 153:29]
  wire [11:0] _T_327; // @[PositDivisionSqrt.scala 153:22]
  wire [14:0] _GEN_11; // @[PositDivisionSqrt.scala 152:93]
  wire [14:0] _T_328; // @[PositDivisionSqrt.scala 152:93]
  wire  _T_330; // @[PositDivisionSqrt.scala 154:33]
  wire  _T_331; // @[PositDivisionSqrt.scala 154:30]
  wire  _T_332; // @[PositDivisionSqrt.scala 154:57]
  wire [14:0] _T_335; // @[Cat.scala 29:58]
  wire [14:0] _T_336; // @[PositDivisionSqrt.scala 154:22]
  wire [14:0] _T_337; // @[PositDivisionSqrt.scala 153:93]
  wire  _T_339; // @[PositDivisionSqrt.scala 155:30]
  wire  _T_340; // @[PositDivisionSqrt.scala 156:83]
  wire [10:0] _T_342; // @[Bitwise.scala 71:12]
  wire [13:0] _GEN_12; // @[PositDivisionSqrt.scala 156:53]
  wire [13:0] _T_343; // @[PositDivisionSqrt.scala 156:53]
  wire [14:0] _GEN_13; // @[PositDivisionSqrt.scala 155:51]
  wire [14:0] _T_344; // @[PositDivisionSqrt.scala 155:51]
  wire [12:0] _T_345; // @[PositDivisionSqrt.scala 157:53]
  wire [14:0] _GEN_14; // @[PositDivisionSqrt.scala 156:89]
  wire [14:0] _T_346; // @[PositDivisionSqrt.scala 156:89]
  wire [14:0] _T_347; // @[PositDivisionSqrt.scala 155:22]
  wire [14:0] trialTerm; // @[PositDivisionSqrt.scala 154:93]
  wire  _T_349; // @[PositDivisionSqrt.scala 162:56]
  wire  _T_350; // @[PositDivisionSqrt.scala 162:40]
  wire [14:0] _T_353; // @[PositDivisionSqrt.scala 163:97]
  wire [14:0] _T_355; // @[PositDivisionSqrt.scala 164:97]
  wire [14:0] _T_356; // @[PositDivisionSqrt.scala 161:92]
  wire [15:0] _T_361; // @[PositDivisionSqrt.scala 168:98]
  wire [14:0] _T_362; // @[PositDivisionSqrt.scala 168:108]
  wire [14:0] _T_364; // @[PositDivisionSqrt.scala 168:112]
  wire [14:0] _T_368; // @[PositDivisionSqrt.scala 169:112]
  wire [14:0] _T_369; // @[PositDivisionSqrt.scala 166:26]
  wire [14:0] trialRem; // @[PositDivisionSqrt.scala 159:27]
  wire  _T_370; // @[PositDivisionSqrt.scala 173:35]
  wire  trIsZero; // @[PositDivisionSqrt.scala 173:25]
  wire  _T_371; // @[PositDivisionSqrt.scala 174:30]
  wire  remIsZero; // @[PositDivisionSqrt.scala 174:25]
  wire  _T_373; // @[PositDivisionSqrt.scala 176:64]
  wire  _T_374; // @[PositDivisionSqrt.scala 176:49]
  wire  _T_375; // @[PositDivisionSqrt.scala 176:29]
  wire  _T_376; // @[PositDivisionSqrt.scala 178:61]
  wire  _T_377; // @[PositDivisionSqrt.scala 178:49]
  wire  _T_379; // @[Mux.scala 87:16]
  wire  newBit; // @[Mux.scala 87:16]
  wire  _T_380; // @[PositDivisionSqrt.scala 183:41]
  wire  _T_381; // @[PositDivisionSqrt.scala 183:51]
  wire  _T_382; // @[PositDivisionSqrt.scala 183:48]
  wire  _T_383; // @[PositDivisionSqrt.scala 183:28]
  wire  _T_386; // @[PositDivisionSqrt.scala 187:39]
  wire  _T_387; // @[PositDivisionSqrt.scala 187:28]
  wire [14:0] _T_390; // @[PositDivisionSqrt.scala 188:47]
  wire [14:0] _T_391; // @[PositDivisionSqrt.scala 188:18]
  wire [12:0] _T_393; // @[PositDivisionSqrt.scala 189:18]
  wire [14:0] _GEN_15; // @[PositDivisionSqrt.scala 188:78]
  wire [14:0] _T_394; // @[PositDivisionSqrt.scala 188:78]
  wire [14:0] _GEN_16; // @[PositDivisionSqrt.scala 190:47]
  wire [14:0] _T_396; // @[PositDivisionSqrt.scala 190:47]
  wire [14:0] _T_397; // @[PositDivisionSqrt.scala 190:18]
  wire [14:0] _T_398; // @[PositDivisionSqrt.scala 189:78]
  wire [1:0] _T_400; // @[PositDivisionSqrt.scala 196:53]
  wire [1:0] sigXBias; // @[PositDivisionSqrt.scala 196:21]
  wire [14:0] _GEN_17; // @[PositDivisionSqrt.scala 197:25]
  wire [14:0] realSigX; // @[PositDivisionSqrt.scala 197:25]
  wire [7:0] _T_403; // @[PositDivisionSqrt.scala 200:97]
  wire [7:0] _T_404; // @[PositDivisionSqrt.scala 201:97]
  wire [7:0] realFrac; // @[PositDivisionSqrt.scala 198:21]
  wire  _T_405; // @[PositDivisionSqrt.scala 205:33]
  wire  _T_406; // @[PositDivisionSqrt.scala 205:58]
  wire  _T_407; // @[PositDivisionSqrt.scala 205:48]
  wire  scaleNeedSub; // @[PositDivisionSqrt.scala 205:23]
  wire  _T_409; // @[PositDivisionSqrt.scala 206:56]
  wire  notNeedSubTwo; // @[PositDivisionSqrt.scala 206:46]
  wire  scaleSubOne; // @[PositDivisionSqrt.scala 207:36]
  wire  _T_410; // @[PositDivisionSqrt.scala 208:38]
  wire  scaleSubTwo; // @[PositDivisionSqrt.scala 208:36]
  wire [1:0] _T_411; // @[Cat.scala 29:58]
  wire [2:0] _T_412; // @[PositDivisionSqrt.scala 209:63]
  wire [6:0] _GEN_18; // @[PositDivisionSqrt.scala 209:31]
  wire [6:0] _T_414; // @[PositDivisionSqrt.scala 209:31]
  wire [6:0] realExp; // @[PositDivisionSqrt.scala 209:31]
  wire  underflow; // @[PositDivisionSqrt.scala 210:31]
  wire  overflow; // @[PositDivisionSqrt.scala 211:31]
  wire  decQ_sign; // @[PositDivisionSqrt.scala 215:33]
  wire [6:0] _T_416; // @[Mux.scala 87:16]
  wire [6:0] _T_417; // @[Mux.scala 87:16]
  wire [2:0] _T_418; // @[PositDivisionSqrt.scala 224:48]
  wire [2:0] _T_419; // @[PositDivisionSqrt.scala 224:64]
  wire [2:0] decQ_grs; // @[PositDivisionSqrt.scala 224:23]
  wire  outValid; // @[PositDivisionSqrt.scala 229:28]
  wire [5:0] _GEN_19; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire [5:0] decQ_scale; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire  _T_425; // @[convert.scala 46:61]
  wire  _T_426; // @[convert.scala 46:52]
  wire  _T_428; // @[convert.scala 46:42]
  wire [4:0] _T_429; // @[convert.scala 48:34]
  wire  _T_430; // @[convert.scala 49:36]
  wire [4:0] _T_432; // @[convert.scala 50:36]
  wire [4:0] _T_433; // @[convert.scala 50:36]
  wire [4:0] _T_434; // @[convert.scala 50:28]
  wire  _T_435; // @[convert.scala 51:31]
  wire  _T_436; // @[convert.scala 52:43]
  wire [13:0] _T_440; // @[Cat.scala 29:58]
  wire [4:0] _T_441; // @[Shift.scala 39:17]
  wire  _T_442; // @[Shift.scala 39:24]
  wire [3:0] _T_443; // @[Shift.scala 40:44]
  wire [5:0] _T_444; // @[Shift.scala 90:30]
  wire [7:0] _T_445; // @[Shift.scala 90:48]
  wire  _T_446; // @[Shift.scala 90:57]
  wire [5:0] _GEN_20; // @[Shift.scala 90:39]
  wire [5:0] _T_447; // @[Shift.scala 90:39]
  wire  _T_448; // @[Shift.scala 12:21]
  wire  _T_449; // @[Shift.scala 12:21]
  wire [7:0] _T_451; // @[Bitwise.scala 71:12]
  wire [13:0] _T_452; // @[Cat.scala 29:58]
  wire [13:0] _T_453; // @[Shift.scala 91:22]
  wire [2:0] _T_454; // @[Shift.scala 92:77]
  wire [9:0] _T_455; // @[Shift.scala 90:30]
  wire [3:0] _T_456; // @[Shift.scala 90:48]
  wire  _T_457; // @[Shift.scala 90:57]
  wire [9:0] _GEN_21; // @[Shift.scala 90:39]
  wire [9:0] _T_458; // @[Shift.scala 90:39]
  wire  _T_459; // @[Shift.scala 12:21]
  wire  _T_460; // @[Shift.scala 12:21]
  wire [3:0] _T_462; // @[Bitwise.scala 71:12]
  wire [13:0] _T_463; // @[Cat.scala 29:58]
  wire [13:0] _T_464; // @[Shift.scala 91:22]
  wire [1:0] _T_465; // @[Shift.scala 92:77]
  wire [11:0] _T_466; // @[Shift.scala 90:30]
  wire [1:0] _T_467; // @[Shift.scala 90:48]
  wire  _T_468; // @[Shift.scala 90:57]
  wire [11:0] _GEN_22; // @[Shift.scala 90:39]
  wire [11:0] _T_469; // @[Shift.scala 90:39]
  wire  _T_470; // @[Shift.scala 12:21]
  wire  _T_471; // @[Shift.scala 12:21]
  wire [1:0] _T_473; // @[Bitwise.scala 71:12]
  wire [13:0] _T_474; // @[Cat.scala 29:58]
  wire [13:0] _T_475; // @[Shift.scala 91:22]
  wire  _T_476; // @[Shift.scala 92:77]
  wire [12:0] _T_477; // @[Shift.scala 90:30]
  wire  _T_478; // @[Shift.scala 90:48]
  wire [12:0] _GEN_23; // @[Shift.scala 90:39]
  wire [12:0] _T_480; // @[Shift.scala 90:39]
  wire  _T_482; // @[Shift.scala 12:21]
  wire [13:0] _T_483; // @[Cat.scala 29:58]
  wire [13:0] _T_484; // @[Shift.scala 91:22]
  wire [13:0] _T_487; // @[Bitwise.scala 71:12]
  wire [13:0] _T_488; // @[Shift.scala 39:10]
  wire  _T_489; // @[convert.scala 55:31]
  wire  _T_490; // @[convert.scala 56:31]
  wire  _T_491; // @[convert.scala 57:31]
  wire  _T_492; // @[convert.scala 58:31]
  wire [10:0] _T_493; // @[convert.scala 59:69]
  wire  _T_494; // @[convert.scala 59:81]
  wire  _T_495; // @[convert.scala 59:50]
  wire  _T_497; // @[convert.scala 60:81]
  wire  _T_498; // @[convert.scala 61:44]
  wire  _T_499; // @[convert.scala 61:52]
  wire  _T_500; // @[convert.scala 61:36]
  wire  _T_501; // @[convert.scala 62:63]
  wire  _T_502; // @[convert.scala 62:103]
  wire  _T_503; // @[convert.scala 62:60]
  wire [10:0] _GEN_24; // @[convert.scala 63:56]
  wire [10:0] _T_506; // @[convert.scala 63:56]
  wire [11:0] _T_507; // @[Cat.scala 29:58]
  wire [11:0] _T_509; // @[Mux.scala 87:16]
  assign _T_1 = io_A[11]; // @[convert.scala 18:24]
  assign _T_2 = io_A[10]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[10:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[9:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[9:2]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[7:4]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8[3:2]; // @[LZD.scala 43:32]
  assign _T_10 = _T_9 != 2'h0; // @[LZD.scala 39:14]
  assign _T_11 = _T_9[1]; // @[LZD.scala 39:21]
  assign _T_12 = _T_9[0]; // @[LZD.scala 39:30]
  assign _T_13 = ~ _T_12; // @[LZD.scala 39:27]
  assign _T_14 = _T_11 | _T_13; // @[LZD.scala 39:25]
  assign _T_15 = {_T_10,_T_14}; // @[Cat.scala 29:58]
  assign _T_16 = _T_8[1:0]; // @[LZD.scala 44:32]
  assign _T_17 = _T_16 != 2'h0; // @[LZD.scala 39:14]
  assign _T_18 = _T_16[1]; // @[LZD.scala 39:21]
  assign _T_19 = _T_16[0]; // @[LZD.scala 39:30]
  assign _T_20 = ~ _T_19; // @[LZD.scala 39:27]
  assign _T_21 = _T_18 | _T_20; // @[LZD.scala 39:25]
  assign _T_22 = {_T_17,_T_21}; // @[Cat.scala 29:58]
  assign _T_23 = _T_15[1]; // @[Shift.scala 12:21]
  assign _T_24 = _T_22[1]; // @[Shift.scala 12:21]
  assign _T_25 = _T_23 | _T_24; // @[LZD.scala 49:16]
  assign _T_26 = ~ _T_24; // @[LZD.scala 49:27]
  assign _T_27 = _T_23 | _T_26; // @[LZD.scala 49:25]
  assign _T_28 = _T_15[0:0]; // @[LZD.scala 49:47]
  assign _T_29 = _T_22[0:0]; // @[LZD.scala 49:59]
  assign _T_30 = _T_23 ? _T_28 : _T_29; // @[LZD.scala 49:35]
  assign _T_32 = {_T_25,_T_27,_T_30}; // @[Cat.scala 29:58]
  assign _T_33 = _T_7[3:0]; // @[LZD.scala 44:32]
  assign _T_34 = _T_33[3:2]; // @[LZD.scala 43:32]
  assign _T_35 = _T_34 != 2'h0; // @[LZD.scala 39:14]
  assign _T_36 = _T_34[1]; // @[LZD.scala 39:21]
  assign _T_37 = _T_34[0]; // @[LZD.scala 39:30]
  assign _T_38 = ~ _T_37; // @[LZD.scala 39:27]
  assign _T_39 = _T_36 | _T_38; // @[LZD.scala 39:25]
  assign _T_40 = {_T_35,_T_39}; // @[Cat.scala 29:58]
  assign _T_41 = _T_33[1:0]; // @[LZD.scala 44:32]
  assign _T_42 = _T_41 != 2'h0; // @[LZD.scala 39:14]
  assign _T_43 = _T_41[1]; // @[LZD.scala 39:21]
  assign _T_44 = _T_41[0]; // @[LZD.scala 39:30]
  assign _T_45 = ~ _T_44; // @[LZD.scala 39:27]
  assign _T_46 = _T_43 | _T_45; // @[LZD.scala 39:25]
  assign _T_47 = {_T_42,_T_46}; // @[Cat.scala 29:58]
  assign _T_48 = _T_40[1]; // @[Shift.scala 12:21]
  assign _T_49 = _T_47[1]; // @[Shift.scala 12:21]
  assign _T_50 = _T_48 | _T_49; // @[LZD.scala 49:16]
  assign _T_51 = ~ _T_49; // @[LZD.scala 49:27]
  assign _T_52 = _T_48 | _T_51; // @[LZD.scala 49:25]
  assign _T_53 = _T_40[0:0]; // @[LZD.scala 49:47]
  assign _T_54 = _T_47[0:0]; // @[LZD.scala 49:59]
  assign _T_55 = _T_48 ? _T_53 : _T_54; // @[LZD.scala 49:35]
  assign _T_57 = {_T_50,_T_52,_T_55}; // @[Cat.scala 29:58]
  assign _T_58 = _T_32[2]; // @[Shift.scala 12:21]
  assign _T_59 = _T_57[2]; // @[Shift.scala 12:21]
  assign _T_60 = _T_58 | _T_59; // @[LZD.scala 49:16]
  assign _T_61 = ~ _T_59; // @[LZD.scala 49:27]
  assign _T_62 = _T_58 | _T_61; // @[LZD.scala 49:25]
  assign _T_63 = _T_32[1:0]; // @[LZD.scala 49:47]
  assign _T_64 = _T_57[1:0]; // @[LZD.scala 49:59]
  assign _T_65 = _T_58 ? _T_63 : _T_64; // @[LZD.scala 49:35]
  assign _T_67 = {_T_60,_T_62,_T_65}; // @[Cat.scala 29:58]
  assign _T_68 = _T_6[1:0]; // @[LZD.scala 44:32]
  assign _T_69 = _T_68 != 2'h0; // @[LZD.scala 39:14]
  assign _T_70 = _T_68[1]; // @[LZD.scala 39:21]
  assign _T_71 = _T_68[0]; // @[LZD.scala 39:30]
  assign _T_72 = ~ _T_71; // @[LZD.scala 39:27]
  assign _T_73 = _T_70 | _T_72; // @[LZD.scala 39:25]
  assign _T_75 = _T_67[3]; // @[Shift.scala 12:21]
  assign _T_77 = {1'h1,_T_69,_T_73}; // @[Cat.scala 29:58]
  assign _T_78 = _T_67[2:0]; // @[LZD.scala 55:32]
  assign _T_79 = _T_75 ? _T_78 : _T_77; // @[LZD.scala 55:20]
  assign _T_80 = {_T_75,_T_79}; // @[Cat.scala 29:58]
  assign _T_81 = ~ _T_80; // @[convert.scala 21:22]
  assign _T_82 = io_A[8:0]; // @[convert.scala 22:36]
  assign _T_83 = _T_81 < 4'h9; // @[Shift.scala 16:24]
  assign _T_85 = _T_81[3]; // @[Shift.scala 12:21]
  assign _T_86 = _T_82[0:0]; // @[Shift.scala 64:52]
  assign _T_88 = {_T_86,8'h0}; // @[Cat.scala 29:58]
  assign _T_89 = _T_85 ? _T_88 : _T_82; // @[Shift.scala 64:27]
  assign _T_90 = _T_81[2:0]; // @[Shift.scala 66:70]
  assign _T_91 = _T_90[2]; // @[Shift.scala 12:21]
  assign _T_92 = _T_89[4:0]; // @[Shift.scala 64:52]
  assign _T_94 = {_T_92,4'h0}; // @[Cat.scala 29:58]
  assign _T_95 = _T_91 ? _T_94 : _T_89; // @[Shift.scala 64:27]
  assign _T_96 = _T_90[1:0]; // @[Shift.scala 66:70]
  assign _T_97 = _T_96[1]; // @[Shift.scala 12:21]
  assign _T_98 = _T_95[6:0]; // @[Shift.scala 64:52]
  assign _T_100 = {_T_98,2'h0}; // @[Cat.scala 29:58]
  assign _T_101 = _T_97 ? _T_100 : _T_95; // @[Shift.scala 64:27]
  assign _T_102 = _T_96[0:0]; // @[Shift.scala 66:70]
  assign _T_104 = _T_101[7:0]; // @[Shift.scala 64:52]
  assign _T_105 = {_T_104,1'h0}; // @[Cat.scala 29:58]
  assign _T_106 = _T_102 ? _T_105 : _T_101; // @[Shift.scala 64:27]
  assign _T_107 = _T_83 ? _T_106 : 9'h0; // @[Shift.scala 16:10]
  assign _T_108 = _T_107[8:8]; // @[convert.scala 23:34]
  assign decA_fraction = _T_107[7:0]; // @[convert.scala 24:34]
  assign _T_110 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_112 = _T_3 ? _T_81 : _T_80; // @[convert.scala 25:42]
  assign _T_115 = ~ _T_108; // @[convert.scala 26:67]
  assign _T_116 = _T_1 ? _T_115 : _T_108; // @[convert.scala 26:51]
  assign _T_117 = {_T_110,_T_112,_T_116}; // @[Cat.scala 29:58]
  assign _T_119 = io_A[10:0]; // @[convert.scala 29:56]
  assign _T_120 = _T_119 != 11'h0; // @[convert.scala 29:60]
  assign _T_121 = ~ _T_120; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_121; // @[convert.scala 29:39]
  assign _T_124 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_124 & _T_121; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_117); // @[convert.scala 32:24]
  assign _T_133 = io_B[11]; // @[convert.scala 18:24]
  assign _T_134 = io_B[10]; // @[convert.scala 18:40]
  assign _T_135 = _T_133 ^ _T_134; // @[convert.scala 18:36]
  assign _T_136 = io_B[10:1]; // @[convert.scala 19:24]
  assign _T_137 = io_B[9:0]; // @[convert.scala 19:43]
  assign _T_138 = _T_136 ^ _T_137; // @[convert.scala 19:39]
  assign _T_139 = _T_138[9:2]; // @[LZD.scala 43:32]
  assign _T_140 = _T_139[7:4]; // @[LZD.scala 43:32]
  assign _T_141 = _T_140[3:2]; // @[LZD.scala 43:32]
  assign _T_142 = _T_141 != 2'h0; // @[LZD.scala 39:14]
  assign _T_143 = _T_141[1]; // @[LZD.scala 39:21]
  assign _T_144 = _T_141[0]; // @[LZD.scala 39:30]
  assign _T_145 = ~ _T_144; // @[LZD.scala 39:27]
  assign _T_146 = _T_143 | _T_145; // @[LZD.scala 39:25]
  assign _T_147 = {_T_142,_T_146}; // @[Cat.scala 29:58]
  assign _T_148 = _T_140[1:0]; // @[LZD.scala 44:32]
  assign _T_149 = _T_148 != 2'h0; // @[LZD.scala 39:14]
  assign _T_150 = _T_148[1]; // @[LZD.scala 39:21]
  assign _T_151 = _T_148[0]; // @[LZD.scala 39:30]
  assign _T_152 = ~ _T_151; // @[LZD.scala 39:27]
  assign _T_153 = _T_150 | _T_152; // @[LZD.scala 39:25]
  assign _T_154 = {_T_149,_T_153}; // @[Cat.scala 29:58]
  assign _T_155 = _T_147[1]; // @[Shift.scala 12:21]
  assign _T_156 = _T_154[1]; // @[Shift.scala 12:21]
  assign _T_157 = _T_155 | _T_156; // @[LZD.scala 49:16]
  assign _T_158 = ~ _T_156; // @[LZD.scala 49:27]
  assign _T_159 = _T_155 | _T_158; // @[LZD.scala 49:25]
  assign _T_160 = _T_147[0:0]; // @[LZD.scala 49:47]
  assign _T_161 = _T_154[0:0]; // @[LZD.scala 49:59]
  assign _T_162 = _T_155 ? _T_160 : _T_161; // @[LZD.scala 49:35]
  assign _T_164 = {_T_157,_T_159,_T_162}; // @[Cat.scala 29:58]
  assign _T_165 = _T_139[3:0]; // @[LZD.scala 44:32]
  assign _T_166 = _T_165[3:2]; // @[LZD.scala 43:32]
  assign _T_167 = _T_166 != 2'h0; // @[LZD.scala 39:14]
  assign _T_168 = _T_166[1]; // @[LZD.scala 39:21]
  assign _T_169 = _T_166[0]; // @[LZD.scala 39:30]
  assign _T_170 = ~ _T_169; // @[LZD.scala 39:27]
  assign _T_171 = _T_168 | _T_170; // @[LZD.scala 39:25]
  assign _T_172 = {_T_167,_T_171}; // @[Cat.scala 29:58]
  assign _T_173 = _T_165[1:0]; // @[LZD.scala 44:32]
  assign _T_174 = _T_173 != 2'h0; // @[LZD.scala 39:14]
  assign _T_175 = _T_173[1]; // @[LZD.scala 39:21]
  assign _T_176 = _T_173[0]; // @[LZD.scala 39:30]
  assign _T_177 = ~ _T_176; // @[LZD.scala 39:27]
  assign _T_178 = _T_175 | _T_177; // @[LZD.scala 39:25]
  assign _T_179 = {_T_174,_T_178}; // @[Cat.scala 29:58]
  assign _T_180 = _T_172[1]; // @[Shift.scala 12:21]
  assign _T_181 = _T_179[1]; // @[Shift.scala 12:21]
  assign _T_182 = _T_180 | _T_181; // @[LZD.scala 49:16]
  assign _T_183 = ~ _T_181; // @[LZD.scala 49:27]
  assign _T_184 = _T_180 | _T_183; // @[LZD.scala 49:25]
  assign _T_185 = _T_172[0:0]; // @[LZD.scala 49:47]
  assign _T_186 = _T_179[0:0]; // @[LZD.scala 49:59]
  assign _T_187 = _T_180 ? _T_185 : _T_186; // @[LZD.scala 49:35]
  assign _T_189 = {_T_182,_T_184,_T_187}; // @[Cat.scala 29:58]
  assign _T_190 = _T_164[2]; // @[Shift.scala 12:21]
  assign _T_191 = _T_189[2]; // @[Shift.scala 12:21]
  assign _T_192 = _T_190 | _T_191; // @[LZD.scala 49:16]
  assign _T_193 = ~ _T_191; // @[LZD.scala 49:27]
  assign _T_194 = _T_190 | _T_193; // @[LZD.scala 49:25]
  assign _T_195 = _T_164[1:0]; // @[LZD.scala 49:47]
  assign _T_196 = _T_189[1:0]; // @[LZD.scala 49:59]
  assign _T_197 = _T_190 ? _T_195 : _T_196; // @[LZD.scala 49:35]
  assign _T_199 = {_T_192,_T_194,_T_197}; // @[Cat.scala 29:58]
  assign _T_200 = _T_138[1:0]; // @[LZD.scala 44:32]
  assign _T_201 = _T_200 != 2'h0; // @[LZD.scala 39:14]
  assign _T_202 = _T_200[1]; // @[LZD.scala 39:21]
  assign _T_203 = _T_200[0]; // @[LZD.scala 39:30]
  assign _T_204 = ~ _T_203; // @[LZD.scala 39:27]
  assign _T_205 = _T_202 | _T_204; // @[LZD.scala 39:25]
  assign _T_207 = _T_199[3]; // @[Shift.scala 12:21]
  assign _T_209 = {1'h1,_T_201,_T_205}; // @[Cat.scala 29:58]
  assign _T_210 = _T_199[2:0]; // @[LZD.scala 55:32]
  assign _T_211 = _T_207 ? _T_210 : _T_209; // @[LZD.scala 55:20]
  assign _T_212 = {_T_207,_T_211}; // @[Cat.scala 29:58]
  assign _T_213 = ~ _T_212; // @[convert.scala 21:22]
  assign _T_214 = io_B[8:0]; // @[convert.scala 22:36]
  assign _T_215 = _T_213 < 4'h9; // @[Shift.scala 16:24]
  assign _T_217 = _T_213[3]; // @[Shift.scala 12:21]
  assign _T_218 = _T_214[0:0]; // @[Shift.scala 64:52]
  assign _T_220 = {_T_218,8'h0}; // @[Cat.scala 29:58]
  assign _T_221 = _T_217 ? _T_220 : _T_214; // @[Shift.scala 64:27]
  assign _T_222 = _T_213[2:0]; // @[Shift.scala 66:70]
  assign _T_223 = _T_222[2]; // @[Shift.scala 12:21]
  assign _T_224 = _T_221[4:0]; // @[Shift.scala 64:52]
  assign _T_226 = {_T_224,4'h0}; // @[Cat.scala 29:58]
  assign _T_227 = _T_223 ? _T_226 : _T_221; // @[Shift.scala 64:27]
  assign _T_228 = _T_222[1:0]; // @[Shift.scala 66:70]
  assign _T_229 = _T_228[1]; // @[Shift.scala 12:21]
  assign _T_230 = _T_227[6:0]; // @[Shift.scala 64:52]
  assign _T_232 = {_T_230,2'h0}; // @[Cat.scala 29:58]
  assign _T_233 = _T_229 ? _T_232 : _T_227; // @[Shift.scala 64:27]
  assign _T_234 = _T_228[0:0]; // @[Shift.scala 66:70]
  assign _T_236 = _T_233[7:0]; // @[Shift.scala 64:52]
  assign _T_237 = {_T_236,1'h0}; // @[Cat.scala 29:58]
  assign _T_238 = _T_234 ? _T_237 : _T_233; // @[Shift.scala 64:27]
  assign _T_239 = _T_215 ? _T_238 : 9'h0; // @[Shift.scala 16:10]
  assign _T_240 = _T_239[8:8]; // @[convert.scala 23:34]
  assign decB_fraction = _T_239[7:0]; // @[convert.scala 24:34]
  assign _T_242 = _T_135 == 1'h0; // @[convert.scala 25:26]
  assign _T_244 = _T_135 ? _T_213 : _T_212; // @[convert.scala 25:42]
  assign _T_247 = ~ _T_240; // @[convert.scala 26:67]
  assign _T_248 = _T_133 ? _T_247 : _T_240; // @[convert.scala 26:51]
  assign _T_249 = {_T_242,_T_244,_T_248}; // @[Cat.scala 29:58]
  assign _T_251 = io_B[10:0]; // @[convert.scala 29:56]
  assign _T_252 = _T_251 != 11'h0; // @[convert.scala 29:60]
  assign _T_253 = ~ _T_252; // @[convert.scala 29:41]
  assign decB_isNaR = _T_133 & _T_253; // @[convert.scala 29:39]
  assign _T_256 = _T_133 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_256 & _T_253; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_249); // @[convert.scala 32:24]
  assign _T_265 = _T_1 ? 3'h7 : 3'h0; // @[Bitwise.scala 71:12]
  assign _T_266 = ~ _T_1; // @[PositDivisionSqrt.scala 80:40]
  assign sigA_S = {_T_265,_T_266,decA_fraction,3'h0}; // @[Cat.scala 29:58]
  assign _T_269 = ~ _T_133; // @[PositDivisionSqrt.scala 82:31]
  assign sigB_S = {_T_133,_T_269,decB_fraction,5'h0}; // @[Cat.scala 29:58]
  assign _T_272 = decA_isNaR == 1'h0; // @[PositDivisionSqrt.scala 85:25]
  assign invalidSqrt = _T_272 & _T_1; // @[PositDivisionSqrt.scala 85:37]
  assign _T_273 = decA_isNaR | invalidSqrt; // @[PositDivisionSqrt.scala 88:42]
  assign _T_274 = decA_isNaR | decB_isNaR; // @[PositDivisionSqrt.scala 89:42]
  assign _T_275 = _T_274 | decB_isZero; // @[PositDivisionSqrt.scala 89:56]
  assign _T_276 = decB_isZero == 1'h0; // @[PositDivisionSqrt.scala 94:46]
  assign _T_277 = decA_isZero & _T_276; // @[PositDivisionSqrt.scala 94:43]
  assign _T_278 = decB_isNaR == 1'h0; // @[PositDivisionSqrt.scala 94:62]
  assign _T_279 = _T_277 & _T_278; // @[PositDivisionSqrt.scala 94:59]
  assign specialCaseA_S = decA_isNaR | decA_isZero; // @[PositDivisionSqrt.scala 97:38]
  assign specialCaseB_S = decB_isNaR | decB_isZero; // @[PositDivisionSqrt.scala 98:38]
  assign _T_280 = specialCaseA_S == 1'h0; // @[PositDivisionSqrt.scala 99:27]
  assign _T_281 = specialCaseB_S == 1'h0; // @[PositDivisionSqrt.scala 99:46]
  assign normalCase_S_div = _T_280 & _T_281; // @[PositDivisionSqrt.scala 99:43]
  assign normalCase_S_sqrt = _T_280 & _T_124; // @[PositDivisionSqrt.scala 100:43]
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div; // @[PositDivisionSqrt.scala 101:30]
  assign sExpQuot_S_div = $signed(decA_scale) - $signed(decB_scale); // @[PositDivisionSqrt.scala 103:38]
  assign _T_284 = decA_scale[0]; // @[PositDivisionSqrt.scala 104:50]
  assign oddSqrt_S = io_sqrtOp & _T_284; // @[PositDivisionSqrt.scala 104:37]
  assign idle = cycleNum == 4'h0; // @[PositDivisionSqrt.scala 109:39]
  assign ready = cycleNum <= 4'h1; // @[PositDivisionSqrt.scala 110:39]
  assign entering = ready & io_inValid; // @[PositDivisionSqrt.scala 111:35]
  assign entering_normalCase = entering & normalCase_S; // @[PositDivisionSqrt.scala 112:38]
  assign _T_285 = sigX_Z[14]; // @[PositDivisionSqrt.scala 113:35]
  assign _T_286 = sigX_Z[12]; // @[PositDivisionSqrt.scala 113:58]
  assign scaleNotChange = _T_285 ^ _T_286; // @[PositDivisionSqrt.scala 113:50]
  assign _T_287 = cycleNum == 4'h3; // @[PositDivisionSqrt.scala 114:39]
  assign skipCycle2 = _T_287 & scaleNotChange; // @[PositDivisionSqrt.scala 114:48]
  assign _T_288 = idle == 1'h0; // @[PositDivisionSqrt.scala 116:8]
  assign _T_289 = _T_288 | io_inValid; // @[PositDivisionSqrt.scala 116:14]
  assign _T_290 = normalCase_S == 1'h0; // @[PositDivisionSqrt.scala 117:32]
  assign _T_291 = entering & _T_290; // @[PositDivisionSqrt.scala 117:30]
  assign _T_293 = io_sqrtOp ? 4'hd : 4'hf; // @[PositDivisionSqrt.scala 119:26]
  assign _T_294 = entering_normalCase ? _T_293 : 4'h0; // @[PositDivisionSqrt.scala 118:20]
  assign _GEN_9 = {{3'd0}, _T_291}; // @[PositDivisionSqrt.scala 117:64]
  assign _T_295 = _GEN_9 | _T_294; // @[PositDivisionSqrt.scala 117:64]
  assign _T_297 = skipCycle2 == 1'h0; // @[PositDivisionSqrt.scala 123:30]
  assign _T_298 = _T_288 & _T_297; // @[PositDivisionSqrt.scala 123:27]
  assign _T_300 = cycleNum - 4'h1; // @[PositDivisionSqrt.scala 123:52]
  assign _T_301 = _T_298 ? _T_300 : 4'h0; // @[PositDivisionSqrt.scala 123:20]
  assign _T_302 = _T_295 | _T_301; // @[PositDivisionSqrt.scala 122:64]
  assign _T_304 = _T_288 & skipCycle2; // @[PositDivisionSqrt.scala 124:27]
  assign _GEN_10 = {{3'd0}, _T_304}; // @[PositDivisionSqrt.scala 123:64]
  assign _T_306 = _T_302 | _GEN_10; // @[PositDivisionSqrt.scala 123:64]
  assign _T_307 = decA_scale[5:1]; // @[PositDivisionSqrt.scala 134:42]
  assign _T_309 = io_sqrtOp == 1'h0; // @[PositDivisionSqrt.scala 137:31]
  assign _T_310 = entering_normalCase & _T_309; // @[PositDivisionSqrt.scala 137:28]
  assign _T_311 = 16'h1 << cycleNum; // @[PositDivisionSqrt.scala 146:22]
  assign bitMask = _T_311[15:2]; // @[PositDivisionSqrt.scala 146:35]
  assign _T_313 = oddSqrt_S == 1'h0; // @[PositDivisionSqrt.scala 148:26]
  assign _T_314 = ready & _T_313; // @[PositDivisionSqrt.scala 148:23]
  assign _T_315 = _T_314 ? sigA_S : 15'h0; // @[PositDivisionSqrt.scala 148:16]
  assign _T_316 = ready & oddSqrt_S; // @[PositDivisionSqrt.scala 149:23]
  assign _T_317 = {sigA_S, 1'h0}; // @[PositDivisionSqrt.scala 149:46]
  assign _T_318 = _T_317[14:0]; // @[PositDivisionSqrt.scala 149:56]
  assign _T_319 = _T_316 ? _T_318 : 15'h0; // @[PositDivisionSqrt.scala 149:16]
  assign _T_320 = _T_315 | _T_319; // @[PositDivisionSqrt.scala 148:66]
  assign _T_321 = ready == 1'h0; // @[PositDivisionSqrt.scala 150:17]
  assign _T_322 = _T_321 ? rem_Z : 15'h0; // @[PositDivisionSqrt.scala 150:16]
  assign rem = _T_320 | _T_322; // @[PositDivisionSqrt.scala 149:66]
  assign _T_324 = ready & _T_309; // @[PositDivisionSqrt.scala 152:29]
  assign _T_325 = _T_324 ? sigB_S : 15'h0; // @[PositDivisionSqrt.scala 152:22]
  assign _T_326 = ready & io_sqrtOp; // @[PositDivisionSqrt.scala 153:29]
  assign _T_327 = _T_326 ? 12'h800 : 12'h0; // @[PositDivisionSqrt.scala 153:22]
  assign _GEN_11 = {{3'd0}, _T_327}; // @[PositDivisionSqrt.scala 152:93]
  assign _T_328 = _T_325 | _GEN_11; // @[PositDivisionSqrt.scala 152:93]
  assign _T_330 = sqrtOp_Z == 1'h0; // @[PositDivisionSqrt.scala 154:33]
  assign _T_331 = _T_321 & _T_330; // @[PositDivisionSqrt.scala 154:30]
  assign _T_332 = ~ signB_Z; // @[PositDivisionSqrt.scala 154:57]
  assign _T_335 = {signB_Z,_T_332,fractB_Z,5'h0}; // @[Cat.scala 29:58]
  assign _T_336 = _T_331 ? _T_335 : 15'h0; // @[PositDivisionSqrt.scala 154:22]
  assign _T_337 = _T_328 | _T_336; // @[PositDivisionSqrt.scala 153:93]
  assign _T_339 = _T_321 & sqrtOp_Z; // @[PositDivisionSqrt.scala 155:30]
  assign _T_340 = rem[14:14]; // @[PositDivisionSqrt.scala 156:83]
  assign _T_342 = _T_340 ? 11'h7ff : 11'h0; // @[Bitwise.scala 71:12]
  assign _GEN_12 = {{3'd0}, _T_342}; // @[PositDivisionSqrt.scala 156:53]
  assign _T_343 = bitMask & _GEN_12; // @[PositDivisionSqrt.scala 156:53]
  assign _GEN_13 = {{1'd0}, _T_343}; // @[PositDivisionSqrt.scala 155:51]
  assign _T_344 = sigX_Z | _GEN_13; // @[PositDivisionSqrt.scala 155:51]
  assign _T_345 = bitMask[13:1]; // @[PositDivisionSqrt.scala 157:53]
  assign _GEN_14 = {{2'd0}, _T_345}; // @[PositDivisionSqrt.scala 156:89]
  assign _T_346 = _T_344 | _GEN_14; // @[PositDivisionSqrt.scala 156:89]
  assign _T_347 = _T_339 ? _T_346 : 15'h0; // @[PositDivisionSqrt.scala 155:22]
  assign trialTerm = _T_337 | _T_347; // @[PositDivisionSqrt.scala 154:93]
  assign _T_349 = trialTerm[14:14]; // @[PositDivisionSqrt.scala 162:56]
  assign _T_350 = _T_340 ^ _T_349; // @[PositDivisionSqrt.scala 162:40]
  assign _T_353 = rem + trialTerm; // @[PositDivisionSqrt.scala 163:97]
  assign _T_355 = rem - trialTerm; // @[PositDivisionSqrt.scala 164:97]
  assign _T_356 = _T_350 ? _T_353 : _T_355; // @[PositDivisionSqrt.scala 161:92]
  assign _T_361 = {rem, 1'h0}; // @[PositDivisionSqrt.scala 168:98]
  assign _T_362 = _T_361[14:0]; // @[PositDivisionSqrt.scala 168:108]
  assign _T_364 = _T_362 + trialTerm; // @[PositDivisionSqrt.scala 168:112]
  assign _T_368 = _T_362 - trialTerm; // @[PositDivisionSqrt.scala 169:112]
  assign _T_369 = _T_350 ? _T_364 : _T_368; // @[PositDivisionSqrt.scala 166:26]
  assign trialRem = ready ? _T_356 : _T_369; // @[PositDivisionSqrt.scala 159:27]
  assign _T_370 = trialRem != 15'h0; // @[PositDivisionSqrt.scala 173:35]
  assign trIsZero = _T_370 == 1'h0; // @[PositDivisionSqrt.scala 173:25]
  assign _T_371 = rem != 15'h0; // @[PositDivisionSqrt.scala 174:30]
  assign remIsZero = _T_371 == 1'h0; // @[PositDivisionSqrt.scala 174:25]
  assign _T_373 = trialRem[14:14]; // @[PositDivisionSqrt.scala 176:64]
  assign _T_374 = _T_349 ^ _T_373; // @[PositDivisionSqrt.scala 176:49]
  assign _T_375 = ~ _T_374; // @[PositDivisionSqrt.scala 176:29]
  assign _T_376 = sigX_Z[14:14]; // @[PositDivisionSqrt.scala 178:61]
  assign _T_377 = ~ _T_376; // @[PositDivisionSqrt.scala 178:49]
  assign _T_379 = remIsZero ? _T_376 : _T_375; // @[Mux.scala 87:16]
  assign newBit = trIsZero ? _T_377 : _T_379; // @[Mux.scala 87:16]
  assign _T_380 = cycleNum > 4'h2; // @[PositDivisionSqrt.scala 183:41]
  assign _T_381 = remIsZero == 1'h0; // @[PositDivisionSqrt.scala 183:51]
  assign _T_382 = _T_380 & _T_381; // @[PositDivisionSqrt.scala 183:48]
  assign _T_383 = entering_normalCase | _T_382; // @[PositDivisionSqrt.scala 183:28]
  assign _T_386 = _T_321 & newBit; // @[PositDivisionSqrt.scala 187:39]
  assign _T_387 = entering_normalCase | _T_386; // @[PositDivisionSqrt.scala 187:28]
  assign _T_390 = {newBit, 14'h0}; // @[PositDivisionSqrt.scala 188:47]
  assign _T_391 = _T_324 ? _T_390 : 15'h0; // @[PositDivisionSqrt.scala 188:18]
  assign _T_393 = _T_326 ? 13'h1000 : 13'h0; // @[PositDivisionSqrt.scala 189:18]
  assign _GEN_15 = {{2'd0}, _T_393}; // @[PositDivisionSqrt.scala 188:78]
  assign _T_394 = _T_391 | _GEN_15; // @[PositDivisionSqrt.scala 188:78]
  assign _GEN_16 = {{1'd0}, bitMask}; // @[PositDivisionSqrt.scala 190:47]
  assign _T_396 = sigX_Z | _GEN_16; // @[PositDivisionSqrt.scala 190:47]
  assign _T_397 = _T_321 ? _T_396 : 15'h0; // @[PositDivisionSqrt.scala 190:18]
  assign _T_398 = _T_394 | _T_397; // @[PositDivisionSqrt.scala 189:78]
  assign _T_400 = {_T_376, 1'h0}; // @[PositDivisionSqrt.scala 196:53]
  assign sigXBias = scaleNotChange ? _T_400 : {{1'd0}, _T_376}; // @[PositDivisionSqrt.scala 196:21]
  assign _GEN_17 = {{13'd0}, sigXBias}; // @[PositDivisionSqrt.scala 197:25]
  assign realSigX = sigX_Z + _GEN_17; // @[PositDivisionSqrt.scala 197:25]
  assign _T_403 = realSigX[11:4]; // @[PositDivisionSqrt.scala 200:97]
  assign _T_404 = realSigX[10:3]; // @[PositDivisionSqrt.scala 201:97]
  assign realFrac = scaleNotChange ? _T_403 : _T_404; // @[PositDivisionSqrt.scala 198:21]
  assign _T_405 = realSigX[14]; // @[PositDivisionSqrt.scala 205:33]
  assign _T_406 = realSigX[12]; // @[PositDivisionSqrt.scala 205:58]
  assign _T_407 = _T_405 ^ _T_406; // @[PositDivisionSqrt.scala 205:48]
  assign scaleNeedSub = ~ _T_407; // @[PositDivisionSqrt.scala 205:23]
  assign _T_409 = realSigX[11]; // @[PositDivisionSqrt.scala 206:56]
  assign notNeedSubTwo = _T_405 ^ _T_409; // @[PositDivisionSqrt.scala 206:46]
  assign scaleSubOne = scaleNeedSub & notNeedSubTwo; // @[PositDivisionSqrt.scala 207:36]
  assign _T_410 = ~ notNeedSubTwo; // @[PositDivisionSqrt.scala 208:38]
  assign scaleSubTwo = scaleNeedSub & _T_410; // @[PositDivisionSqrt.scala 208:36]
  assign _T_411 = {scaleSubTwo,scaleSubOne}; // @[Cat.scala 29:58]
  assign _T_412 = {1'b0,$signed(_T_411)}; // @[PositDivisionSqrt.scala 209:63]
  assign _GEN_18 = {{4{_T_412[2]}},_T_412}; // @[PositDivisionSqrt.scala 209:31]
  assign _T_414 = $signed(scale_Z) - $signed(_GEN_18); // @[PositDivisionSqrt.scala 209:31]
  assign realExp = $signed(_T_414); // @[PositDivisionSqrt.scala 209:31]
  assign underflow = $signed(realExp) < $signed(-7'sh15); // @[PositDivisionSqrt.scala 210:31]
  assign overflow = $signed(realExp) > $signed(7'sh14); // @[PositDivisionSqrt.scala 211:31]
  assign decQ_sign = realSigX[14:14]; // @[PositDivisionSqrt.scala 215:33]
  assign _T_416 = underflow ? $signed(-7'sh15) : $signed(realExp); // @[Mux.scala 87:16]
  assign _T_417 = overflow ? $signed(7'sh14) : $signed(_T_416); // @[Mux.scala 87:16]
  assign _T_418 = realSigX[3:1]; // @[PositDivisionSqrt.scala 224:48]
  assign _T_419 = realSigX[2:0]; // @[PositDivisionSqrt.scala 224:64]
  assign decQ_grs = scaleNotChange ? _T_418 : _T_419; // @[PositDivisionSqrt.scala 224:23]
  assign outValid = cycleNum == 4'h1; // @[PositDivisionSqrt.scala 229:28]
  assign _GEN_19 = _T_417[5:0]; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign decQ_scale = $signed(_GEN_19); // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign _T_425 = decQ_scale[0]; // @[convert.scala 46:61]
  assign _T_426 = ~ _T_425; // @[convert.scala 46:52]
  assign _T_428 = decQ_sign ? _T_426 : _T_425; // @[convert.scala 46:42]
  assign _T_429 = decQ_scale[5:1]; // @[convert.scala 48:34]
  assign _T_430 = _T_429[4:4]; // @[convert.scala 49:36]
  assign _T_432 = ~ _T_429; // @[convert.scala 50:36]
  assign _T_433 = $signed(_T_432); // @[convert.scala 50:36]
  assign _T_434 = _T_430 ? $signed(_T_433) : $signed(_T_429); // @[convert.scala 50:28]
  assign _T_435 = _T_430 ^ decQ_sign; // @[convert.scala 51:31]
  assign _T_436 = ~ _T_435; // @[convert.scala 52:43]
  assign _T_440 = {_T_436,_T_435,_T_428,realFrac,decQ_grs}; // @[Cat.scala 29:58]
  assign _T_441 = $unsigned(_T_434); // @[Shift.scala 39:17]
  assign _T_442 = _T_441 < 5'he; // @[Shift.scala 39:24]
  assign _T_443 = _T_434[3:0]; // @[Shift.scala 40:44]
  assign _T_444 = _T_440[13:8]; // @[Shift.scala 90:30]
  assign _T_445 = _T_440[7:0]; // @[Shift.scala 90:48]
  assign _T_446 = _T_445 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_20 = {{5'd0}, _T_446}; // @[Shift.scala 90:39]
  assign _T_447 = _T_444 | _GEN_20; // @[Shift.scala 90:39]
  assign _T_448 = _T_443[3]; // @[Shift.scala 12:21]
  assign _T_449 = _T_440[13]; // @[Shift.scala 12:21]
  assign _T_451 = _T_449 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_452 = {_T_451,_T_447}; // @[Cat.scala 29:58]
  assign _T_453 = _T_448 ? _T_452 : _T_440; // @[Shift.scala 91:22]
  assign _T_454 = _T_443[2:0]; // @[Shift.scala 92:77]
  assign _T_455 = _T_453[13:4]; // @[Shift.scala 90:30]
  assign _T_456 = _T_453[3:0]; // @[Shift.scala 90:48]
  assign _T_457 = _T_456 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_21 = {{9'd0}, _T_457}; // @[Shift.scala 90:39]
  assign _T_458 = _T_455 | _GEN_21; // @[Shift.scala 90:39]
  assign _T_459 = _T_454[2]; // @[Shift.scala 12:21]
  assign _T_460 = _T_453[13]; // @[Shift.scala 12:21]
  assign _T_462 = _T_460 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_463 = {_T_462,_T_458}; // @[Cat.scala 29:58]
  assign _T_464 = _T_459 ? _T_463 : _T_453; // @[Shift.scala 91:22]
  assign _T_465 = _T_454[1:0]; // @[Shift.scala 92:77]
  assign _T_466 = _T_464[13:2]; // @[Shift.scala 90:30]
  assign _T_467 = _T_464[1:0]; // @[Shift.scala 90:48]
  assign _T_468 = _T_467 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_22 = {{11'd0}, _T_468}; // @[Shift.scala 90:39]
  assign _T_469 = _T_466 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_470 = _T_465[1]; // @[Shift.scala 12:21]
  assign _T_471 = _T_464[13]; // @[Shift.scala 12:21]
  assign _T_473 = _T_471 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_474 = {_T_473,_T_469}; // @[Cat.scala 29:58]
  assign _T_475 = _T_470 ? _T_474 : _T_464; // @[Shift.scala 91:22]
  assign _T_476 = _T_465[0:0]; // @[Shift.scala 92:77]
  assign _T_477 = _T_475[13:1]; // @[Shift.scala 90:30]
  assign _T_478 = _T_475[0:0]; // @[Shift.scala 90:48]
  assign _GEN_23 = {{12'd0}, _T_478}; // @[Shift.scala 90:39]
  assign _T_480 = _T_477 | _GEN_23; // @[Shift.scala 90:39]
  assign _T_482 = _T_475[13]; // @[Shift.scala 12:21]
  assign _T_483 = {_T_482,_T_480}; // @[Cat.scala 29:58]
  assign _T_484 = _T_476 ? _T_483 : _T_475; // @[Shift.scala 91:22]
  assign _T_487 = _T_449 ? 14'h3fff : 14'h0; // @[Bitwise.scala 71:12]
  assign _T_488 = _T_442 ? _T_484 : _T_487; // @[Shift.scala 39:10]
  assign _T_489 = _T_488[3]; // @[convert.scala 55:31]
  assign _T_490 = _T_488[2]; // @[convert.scala 56:31]
  assign _T_491 = _T_488[1]; // @[convert.scala 57:31]
  assign _T_492 = _T_488[0]; // @[convert.scala 58:31]
  assign _T_493 = _T_488[13:3]; // @[convert.scala 59:69]
  assign _T_494 = _T_493 != 11'h0; // @[convert.scala 59:81]
  assign _T_495 = ~ _T_494; // @[convert.scala 59:50]
  assign _T_497 = _T_493 == 11'h7ff; // @[convert.scala 60:81]
  assign _T_498 = _T_489 | _T_491; // @[convert.scala 61:44]
  assign _T_499 = _T_498 | _T_492; // @[convert.scala 61:52]
  assign _T_500 = _T_490 & _T_499; // @[convert.scala 61:36]
  assign _T_501 = ~ _T_497; // @[convert.scala 62:63]
  assign _T_502 = _T_501 & _T_500; // @[convert.scala 62:103]
  assign _T_503 = _T_495 | _T_502; // @[convert.scala 62:60]
  assign _GEN_24 = {{10'd0}, _T_503}; // @[convert.scala 63:56]
  assign _T_506 = _T_493 + _GEN_24; // @[convert.scala 63:56]
  assign _T_507 = {decQ_sign,_T_506}; // @[Cat.scala 29:58]
  assign _T_509 = isZero_Z ? 12'h0 : _T_507; // @[Mux.scala 87:16]
  assign io_inReady = cycleNum <= 4'h1; // @[PositDivisionSqrt.scala 231:17]
  assign io_diviValid = outValid & _T_330; // @[PositDivisionSqrt.scala 232:17]
  assign io_sqrtValid = outValid & sqrtOp_Z; // @[PositDivisionSqrt.scala 233:17]
  assign io_invalidExc = isNaR_Z; // @[PositDivisionSqrt.scala 234:17]
  assign io_Q = isNaR_Z ? 12'h800 : _T_509; // @[PositDivisionSqrt.scala 235:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleNum = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sqrtOp_Z = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  isNaR_Z = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  isZero_Z = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  scale_Z = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  signB_Z = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fractB_Z = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rem_Z = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sigX_Z = _RAND_8[14:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      cycleNum <= 4'h0;
    end else begin
      if (_T_289) begin
        cycleNum <= _T_306;
      end
    end
    if (entering) begin
      sqrtOp_Z <= io_sqrtOp;
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isNaR_Z <= _T_273;
      end else begin
        isNaR_Z <= _T_275;
      end
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isZero_Z <= decA_isZero;
      end else begin
        isZero_Z <= _T_279;
      end
    end
    if (entering_normalCase) begin
      if (io_sqrtOp) begin
        scale_Z <= {{2{_T_307[4]}},_T_307};
      end else begin
        scale_Z <= sExpQuot_S_div;
      end
    end
    if (_T_310) begin
      signB_Z <= _T_133;
    end
    if (_T_310) begin
      fractB_Z <= decB_fraction;
    end
    if (_T_383) begin
      if (ready) begin
        if (_T_350) begin
          rem_Z <= _T_353;
        end else begin
          rem_Z <= _T_355;
        end
      end else begin
        if (_T_350) begin
          rem_Z <= _T_364;
        end else begin
          rem_Z <= _T_368;
        end
      end
    end
    if (_T_387) begin
      sigX_Z <= _T_398;
    end
  end
endmodule
