module PositDivSqrter32_1(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input  [31:0] io_A,
  input  [31:0] io_B,
  output        io_diviValid,
  output        io_sqrtValid,
  output        io_invalidExc,
  output [31:0] io_Q
);
  reg [5:0] cycleNum; // @[PositDivisionSqrt.scala 63:26]
  reg [31:0] _RAND_0;
  reg  sqrtOp_Z; // @[PositDivisionSqrt.scala 65:22]
  reg [31:0] _RAND_1;
  reg  isNaR_Z; // @[PositDivisionSqrt.scala 66:22]
  reg [31:0] _RAND_2;
  reg  isZero_Z; // @[PositDivisionSqrt.scala 67:22]
  reg [31:0] _RAND_3;
  reg [7:0] scale_Z; // @[PositDivisionSqrt.scala 68:22]
  reg [31:0] _RAND_4;
  reg  signB_Z; // @[PositDivisionSqrt.scala 69:28]
  reg [31:0] _RAND_5;
  reg [27:0] fractB_Z; // @[PositDivisionSqrt.scala 70:22]
  reg [31:0] _RAND_6;
  reg [34:0] rem_Z; // @[PositDivisionSqrt.scala 71:22]
  reg [63:0] _RAND_7;
  reg [34:0] sigX_Z; // @[PositDivisionSqrt.scala 72:22]
  reg [63:0] _RAND_8;
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [29:0] _T_4; // @[convert.scala 19:24]
  wire [29:0] _T_5; // @[convert.scala 19:43]
  wire [29:0] _T_6; // @[convert.scala 19:39]
  wire [15:0] _T_7; // @[LZD.scala 43:32]
  wire [7:0] _T_8; // @[LZD.scala 43:32]
  wire [3:0] _T_9; // @[LZD.scala 43:32]
  wire [1:0] _T_10; // @[LZD.scala 43:32]
  wire  _T_11; // @[LZD.scala 39:14]
  wire  _T_12; // @[LZD.scala 39:21]
  wire  _T_13; // @[LZD.scala 39:30]
  wire  _T_14; // @[LZD.scala 39:27]
  wire  _T_15; // @[LZD.scala 39:25]
  wire [1:0] _T_16; // @[Cat.scala 29:58]
  wire [1:0] _T_17; // @[LZD.scala 44:32]
  wire  _T_18; // @[LZD.scala 39:14]
  wire  _T_19; // @[LZD.scala 39:21]
  wire  _T_20; // @[LZD.scala 39:30]
  wire  _T_21; // @[LZD.scala 39:27]
  wire  _T_22; // @[LZD.scala 39:25]
  wire [1:0] _T_23; // @[Cat.scala 29:58]
  wire  _T_24; // @[Shift.scala 12:21]
  wire  _T_25; // @[Shift.scala 12:21]
  wire  _T_26; // @[LZD.scala 49:16]
  wire  _T_27; // @[LZD.scala 49:27]
  wire  _T_28; // @[LZD.scala 49:25]
  wire  _T_29; // @[LZD.scala 49:47]
  wire  _T_30; // @[LZD.scala 49:59]
  wire  _T_31; // @[LZD.scala 49:35]
  wire [2:0] _T_33; // @[Cat.scala 29:58]
  wire [3:0] _T_34; // @[LZD.scala 44:32]
  wire [1:0] _T_35; // @[LZD.scala 43:32]
  wire  _T_36; // @[LZD.scala 39:14]
  wire  _T_37; // @[LZD.scala 39:21]
  wire  _T_38; // @[LZD.scala 39:30]
  wire  _T_39; // @[LZD.scala 39:27]
  wire  _T_40; // @[LZD.scala 39:25]
  wire [1:0] _T_41; // @[Cat.scala 29:58]
  wire [1:0] _T_42; // @[LZD.scala 44:32]
  wire  _T_43; // @[LZD.scala 39:14]
  wire  _T_44; // @[LZD.scala 39:21]
  wire  _T_45; // @[LZD.scala 39:30]
  wire  _T_46; // @[LZD.scala 39:27]
  wire  _T_47; // @[LZD.scala 39:25]
  wire [1:0] _T_48; // @[Cat.scala 29:58]
  wire  _T_49; // @[Shift.scala 12:21]
  wire  _T_50; // @[Shift.scala 12:21]
  wire  _T_51; // @[LZD.scala 49:16]
  wire  _T_52; // @[LZD.scala 49:27]
  wire  _T_53; // @[LZD.scala 49:25]
  wire  _T_54; // @[LZD.scala 49:47]
  wire  _T_55; // @[LZD.scala 49:59]
  wire  _T_56; // @[LZD.scala 49:35]
  wire [2:0] _T_58; // @[Cat.scala 29:58]
  wire  _T_59; // @[Shift.scala 12:21]
  wire  _T_60; // @[Shift.scala 12:21]
  wire  _T_61; // @[LZD.scala 49:16]
  wire  _T_62; // @[LZD.scala 49:27]
  wire  _T_63; // @[LZD.scala 49:25]
  wire [1:0] _T_64; // @[LZD.scala 49:47]
  wire [1:0] _T_65; // @[LZD.scala 49:59]
  wire [1:0] _T_66; // @[LZD.scala 49:35]
  wire [3:0] _T_68; // @[Cat.scala 29:58]
  wire [7:0] _T_69; // @[LZD.scala 44:32]
  wire [3:0] _T_70; // @[LZD.scala 43:32]
  wire [1:0] _T_71; // @[LZD.scala 43:32]
  wire  _T_72; // @[LZD.scala 39:14]
  wire  _T_73; // @[LZD.scala 39:21]
  wire  _T_74; // @[LZD.scala 39:30]
  wire  _T_75; // @[LZD.scala 39:27]
  wire  _T_76; // @[LZD.scala 39:25]
  wire [1:0] _T_77; // @[Cat.scala 29:58]
  wire [1:0] _T_78; // @[LZD.scala 44:32]
  wire  _T_79; // @[LZD.scala 39:14]
  wire  _T_80; // @[LZD.scala 39:21]
  wire  _T_81; // @[LZD.scala 39:30]
  wire  _T_82; // @[LZD.scala 39:27]
  wire  _T_83; // @[LZD.scala 39:25]
  wire [1:0] _T_84; // @[Cat.scala 29:58]
  wire  _T_85; // @[Shift.scala 12:21]
  wire  _T_86; // @[Shift.scala 12:21]
  wire  _T_87; // @[LZD.scala 49:16]
  wire  _T_88; // @[LZD.scala 49:27]
  wire  _T_89; // @[LZD.scala 49:25]
  wire  _T_90; // @[LZD.scala 49:47]
  wire  _T_91; // @[LZD.scala 49:59]
  wire  _T_92; // @[LZD.scala 49:35]
  wire [2:0] _T_94; // @[Cat.scala 29:58]
  wire [3:0] _T_95; // @[LZD.scala 44:32]
  wire [1:0] _T_96; // @[LZD.scala 43:32]
  wire  _T_97; // @[LZD.scala 39:14]
  wire  _T_98; // @[LZD.scala 39:21]
  wire  _T_99; // @[LZD.scala 39:30]
  wire  _T_100; // @[LZD.scala 39:27]
  wire  _T_101; // @[LZD.scala 39:25]
  wire [1:0] _T_102; // @[Cat.scala 29:58]
  wire [1:0] _T_103; // @[LZD.scala 44:32]
  wire  _T_104; // @[LZD.scala 39:14]
  wire  _T_105; // @[LZD.scala 39:21]
  wire  _T_106; // @[LZD.scala 39:30]
  wire  _T_107; // @[LZD.scala 39:27]
  wire  _T_108; // @[LZD.scala 39:25]
  wire [1:0] _T_109; // @[Cat.scala 29:58]
  wire  _T_110; // @[Shift.scala 12:21]
  wire  _T_111; // @[Shift.scala 12:21]
  wire  _T_112; // @[LZD.scala 49:16]
  wire  _T_113; // @[LZD.scala 49:27]
  wire  _T_114; // @[LZD.scala 49:25]
  wire  _T_115; // @[LZD.scala 49:47]
  wire  _T_116; // @[LZD.scala 49:59]
  wire  _T_117; // @[LZD.scala 49:35]
  wire [2:0] _T_119; // @[Cat.scala 29:58]
  wire  _T_120; // @[Shift.scala 12:21]
  wire  _T_121; // @[Shift.scala 12:21]
  wire  _T_122; // @[LZD.scala 49:16]
  wire  _T_123; // @[LZD.scala 49:27]
  wire  _T_124; // @[LZD.scala 49:25]
  wire [1:0] _T_125; // @[LZD.scala 49:47]
  wire [1:0] _T_126; // @[LZD.scala 49:59]
  wire [1:0] _T_127; // @[LZD.scala 49:35]
  wire [3:0] _T_129; // @[Cat.scala 29:58]
  wire  _T_130; // @[Shift.scala 12:21]
  wire  _T_131; // @[Shift.scala 12:21]
  wire  _T_132; // @[LZD.scala 49:16]
  wire  _T_133; // @[LZD.scala 49:27]
  wire  _T_134; // @[LZD.scala 49:25]
  wire [2:0] _T_135; // @[LZD.scala 49:47]
  wire [2:0] _T_136; // @[LZD.scala 49:59]
  wire [2:0] _T_137; // @[LZD.scala 49:35]
  wire [4:0] _T_139; // @[Cat.scala 29:58]
  wire [13:0] _T_140; // @[LZD.scala 44:32]
  wire [7:0] _T_141; // @[LZD.scala 43:32]
  wire [3:0] _T_142; // @[LZD.scala 43:32]
  wire [1:0] _T_143; // @[LZD.scala 43:32]
  wire  _T_144; // @[LZD.scala 39:14]
  wire  _T_145; // @[LZD.scala 39:21]
  wire  _T_146; // @[LZD.scala 39:30]
  wire  _T_147; // @[LZD.scala 39:27]
  wire  _T_148; // @[LZD.scala 39:25]
  wire [1:0] _T_149; // @[Cat.scala 29:58]
  wire [1:0] _T_150; // @[LZD.scala 44:32]
  wire  _T_151; // @[LZD.scala 39:14]
  wire  _T_152; // @[LZD.scala 39:21]
  wire  _T_153; // @[LZD.scala 39:30]
  wire  _T_154; // @[LZD.scala 39:27]
  wire  _T_155; // @[LZD.scala 39:25]
  wire [1:0] _T_156; // @[Cat.scala 29:58]
  wire  _T_157; // @[Shift.scala 12:21]
  wire  _T_158; // @[Shift.scala 12:21]
  wire  _T_159; // @[LZD.scala 49:16]
  wire  _T_160; // @[LZD.scala 49:27]
  wire  _T_161; // @[LZD.scala 49:25]
  wire  _T_162; // @[LZD.scala 49:47]
  wire  _T_163; // @[LZD.scala 49:59]
  wire  _T_164; // @[LZD.scala 49:35]
  wire [2:0] _T_166; // @[Cat.scala 29:58]
  wire [3:0] _T_167; // @[LZD.scala 44:32]
  wire [1:0] _T_168; // @[LZD.scala 43:32]
  wire  _T_169; // @[LZD.scala 39:14]
  wire  _T_170; // @[LZD.scala 39:21]
  wire  _T_171; // @[LZD.scala 39:30]
  wire  _T_172; // @[LZD.scala 39:27]
  wire  _T_173; // @[LZD.scala 39:25]
  wire [1:0] _T_174; // @[Cat.scala 29:58]
  wire [1:0] _T_175; // @[LZD.scala 44:32]
  wire  _T_176; // @[LZD.scala 39:14]
  wire  _T_177; // @[LZD.scala 39:21]
  wire  _T_178; // @[LZD.scala 39:30]
  wire  _T_179; // @[LZD.scala 39:27]
  wire  _T_180; // @[LZD.scala 39:25]
  wire [1:0] _T_181; // @[Cat.scala 29:58]
  wire  _T_182; // @[Shift.scala 12:21]
  wire  _T_183; // @[Shift.scala 12:21]
  wire  _T_184; // @[LZD.scala 49:16]
  wire  _T_185; // @[LZD.scala 49:27]
  wire  _T_186; // @[LZD.scala 49:25]
  wire  _T_187; // @[LZD.scala 49:47]
  wire  _T_188; // @[LZD.scala 49:59]
  wire  _T_189; // @[LZD.scala 49:35]
  wire [2:0] _T_191; // @[Cat.scala 29:58]
  wire  _T_192; // @[Shift.scala 12:21]
  wire  _T_193; // @[Shift.scala 12:21]
  wire  _T_194; // @[LZD.scala 49:16]
  wire  _T_195; // @[LZD.scala 49:27]
  wire  _T_196; // @[LZD.scala 49:25]
  wire [1:0] _T_197; // @[LZD.scala 49:47]
  wire [1:0] _T_198; // @[LZD.scala 49:59]
  wire [1:0] _T_199; // @[LZD.scala 49:35]
  wire [3:0] _T_201; // @[Cat.scala 29:58]
  wire [5:0] _T_202; // @[LZD.scala 44:32]
  wire [3:0] _T_203; // @[LZD.scala 43:32]
  wire [1:0] _T_204; // @[LZD.scala 43:32]
  wire  _T_205; // @[LZD.scala 39:14]
  wire  _T_206; // @[LZD.scala 39:21]
  wire  _T_207; // @[LZD.scala 39:30]
  wire  _T_208; // @[LZD.scala 39:27]
  wire  _T_209; // @[LZD.scala 39:25]
  wire [1:0] _T_210; // @[Cat.scala 29:58]
  wire [1:0] _T_211; // @[LZD.scala 44:32]
  wire  _T_212; // @[LZD.scala 39:14]
  wire  _T_213; // @[LZD.scala 39:21]
  wire  _T_214; // @[LZD.scala 39:30]
  wire  _T_215; // @[LZD.scala 39:27]
  wire  _T_216; // @[LZD.scala 39:25]
  wire [1:0] _T_217; // @[Cat.scala 29:58]
  wire  _T_218; // @[Shift.scala 12:21]
  wire  _T_219; // @[Shift.scala 12:21]
  wire  _T_220; // @[LZD.scala 49:16]
  wire  _T_221; // @[LZD.scala 49:27]
  wire  _T_222; // @[LZD.scala 49:25]
  wire  _T_223; // @[LZD.scala 49:47]
  wire  _T_224; // @[LZD.scala 49:59]
  wire  _T_225; // @[LZD.scala 49:35]
  wire [2:0] _T_227; // @[Cat.scala 29:58]
  wire [1:0] _T_228; // @[LZD.scala 44:32]
  wire  _T_229; // @[LZD.scala 39:14]
  wire  _T_230; // @[LZD.scala 39:21]
  wire  _T_231; // @[LZD.scala 39:30]
  wire  _T_232; // @[LZD.scala 39:27]
  wire  _T_233; // @[LZD.scala 39:25]
  wire [1:0] _T_234; // @[Cat.scala 29:58]
  wire  _T_235; // @[Shift.scala 12:21]
  wire [1:0] _T_237; // @[LZD.scala 55:32]
  wire [1:0] _T_238; // @[LZD.scala 55:20]
  wire [2:0] _T_239; // @[Cat.scala 29:58]
  wire  _T_240; // @[Shift.scala 12:21]
  wire [2:0] _T_242; // @[LZD.scala 55:32]
  wire [2:0] _T_243; // @[LZD.scala 55:20]
  wire [3:0] _T_244; // @[Cat.scala 29:58]
  wire  _T_245; // @[Shift.scala 12:21]
  wire [3:0] _T_247; // @[LZD.scala 55:32]
  wire [3:0] _T_248; // @[LZD.scala 55:20]
  wire [4:0] _T_249; // @[Cat.scala 29:58]
  wire [4:0] _T_250; // @[convert.scala 21:22]
  wire [28:0] _T_251; // @[convert.scala 22:36]
  wire  _T_252; // @[Shift.scala 16:24]
  wire  _T_254; // @[Shift.scala 12:21]
  wire [12:0] _T_255; // @[Shift.scala 64:52]
  wire [28:0] _T_257; // @[Cat.scala 29:58]
  wire [28:0] _T_258; // @[Shift.scala 64:27]
  wire [3:0] _T_259; // @[Shift.scala 66:70]
  wire  _T_260; // @[Shift.scala 12:21]
  wire [20:0] _T_261; // @[Shift.scala 64:52]
  wire [28:0] _T_263; // @[Cat.scala 29:58]
  wire [28:0] _T_264; // @[Shift.scala 64:27]
  wire [2:0] _T_265; // @[Shift.scala 66:70]
  wire  _T_266; // @[Shift.scala 12:21]
  wire [24:0] _T_267; // @[Shift.scala 64:52]
  wire [28:0] _T_269; // @[Cat.scala 29:58]
  wire [28:0] _T_270; // @[Shift.scala 64:27]
  wire [1:0] _T_271; // @[Shift.scala 66:70]
  wire  _T_272; // @[Shift.scala 12:21]
  wire [26:0] _T_273; // @[Shift.scala 64:52]
  wire [28:0] _T_275; // @[Cat.scala 29:58]
  wire [28:0] _T_276; // @[Shift.scala 64:27]
  wire  _T_277; // @[Shift.scala 66:70]
  wire [27:0] _T_279; // @[Shift.scala 64:52]
  wire [28:0] _T_280; // @[Cat.scala 29:58]
  wire [28:0] _T_281; // @[Shift.scala 64:27]
  wire [28:0] _T_282; // @[Shift.scala 16:10]
  wire  _T_283; // @[convert.scala 23:34]
  wire [27:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_285; // @[convert.scala 25:26]
  wire [4:0] _T_287; // @[convert.scala 25:42]
  wire  _T_290; // @[convert.scala 26:67]
  wire  _T_291; // @[convert.scala 26:51]
  wire [6:0] _T_292; // @[Cat.scala 29:58]
  wire [30:0] _T_294; // @[convert.scala 29:56]
  wire  _T_295; // @[convert.scala 29:60]
  wire  _T_296; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_299; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [6:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_308; // @[convert.scala 18:24]
  wire  _T_309; // @[convert.scala 18:40]
  wire  _T_310; // @[convert.scala 18:36]
  wire [29:0] _T_311; // @[convert.scala 19:24]
  wire [29:0] _T_312; // @[convert.scala 19:43]
  wire [29:0] _T_313; // @[convert.scala 19:39]
  wire [15:0] _T_314; // @[LZD.scala 43:32]
  wire [7:0] _T_315; // @[LZD.scala 43:32]
  wire [3:0] _T_316; // @[LZD.scala 43:32]
  wire [1:0] _T_317; // @[LZD.scala 43:32]
  wire  _T_318; // @[LZD.scala 39:14]
  wire  _T_319; // @[LZD.scala 39:21]
  wire  _T_320; // @[LZD.scala 39:30]
  wire  _T_321; // @[LZD.scala 39:27]
  wire  _T_322; // @[LZD.scala 39:25]
  wire [1:0] _T_323; // @[Cat.scala 29:58]
  wire [1:0] _T_324; // @[LZD.scala 44:32]
  wire  _T_325; // @[LZD.scala 39:14]
  wire  _T_326; // @[LZD.scala 39:21]
  wire  _T_327; // @[LZD.scala 39:30]
  wire  _T_328; // @[LZD.scala 39:27]
  wire  _T_329; // @[LZD.scala 39:25]
  wire [1:0] _T_330; // @[Cat.scala 29:58]
  wire  _T_331; // @[Shift.scala 12:21]
  wire  _T_332; // @[Shift.scala 12:21]
  wire  _T_333; // @[LZD.scala 49:16]
  wire  _T_334; // @[LZD.scala 49:27]
  wire  _T_335; // @[LZD.scala 49:25]
  wire  _T_336; // @[LZD.scala 49:47]
  wire  _T_337; // @[LZD.scala 49:59]
  wire  _T_338; // @[LZD.scala 49:35]
  wire [2:0] _T_340; // @[Cat.scala 29:58]
  wire [3:0] _T_341; // @[LZD.scala 44:32]
  wire [1:0] _T_342; // @[LZD.scala 43:32]
  wire  _T_343; // @[LZD.scala 39:14]
  wire  _T_344; // @[LZD.scala 39:21]
  wire  _T_345; // @[LZD.scala 39:30]
  wire  _T_346; // @[LZD.scala 39:27]
  wire  _T_347; // @[LZD.scala 39:25]
  wire [1:0] _T_348; // @[Cat.scala 29:58]
  wire [1:0] _T_349; // @[LZD.scala 44:32]
  wire  _T_350; // @[LZD.scala 39:14]
  wire  _T_351; // @[LZD.scala 39:21]
  wire  _T_352; // @[LZD.scala 39:30]
  wire  _T_353; // @[LZD.scala 39:27]
  wire  _T_354; // @[LZD.scala 39:25]
  wire [1:0] _T_355; // @[Cat.scala 29:58]
  wire  _T_356; // @[Shift.scala 12:21]
  wire  _T_357; // @[Shift.scala 12:21]
  wire  _T_358; // @[LZD.scala 49:16]
  wire  _T_359; // @[LZD.scala 49:27]
  wire  _T_360; // @[LZD.scala 49:25]
  wire  _T_361; // @[LZD.scala 49:47]
  wire  _T_362; // @[LZD.scala 49:59]
  wire  _T_363; // @[LZD.scala 49:35]
  wire [2:0] _T_365; // @[Cat.scala 29:58]
  wire  _T_366; // @[Shift.scala 12:21]
  wire  _T_367; // @[Shift.scala 12:21]
  wire  _T_368; // @[LZD.scala 49:16]
  wire  _T_369; // @[LZD.scala 49:27]
  wire  _T_370; // @[LZD.scala 49:25]
  wire [1:0] _T_371; // @[LZD.scala 49:47]
  wire [1:0] _T_372; // @[LZD.scala 49:59]
  wire [1:0] _T_373; // @[LZD.scala 49:35]
  wire [3:0] _T_375; // @[Cat.scala 29:58]
  wire [7:0] _T_376; // @[LZD.scala 44:32]
  wire [3:0] _T_377; // @[LZD.scala 43:32]
  wire [1:0] _T_378; // @[LZD.scala 43:32]
  wire  _T_379; // @[LZD.scala 39:14]
  wire  _T_380; // @[LZD.scala 39:21]
  wire  _T_381; // @[LZD.scala 39:30]
  wire  _T_382; // @[LZD.scala 39:27]
  wire  _T_383; // @[LZD.scala 39:25]
  wire [1:0] _T_384; // @[Cat.scala 29:58]
  wire [1:0] _T_385; // @[LZD.scala 44:32]
  wire  _T_386; // @[LZD.scala 39:14]
  wire  _T_387; // @[LZD.scala 39:21]
  wire  _T_388; // @[LZD.scala 39:30]
  wire  _T_389; // @[LZD.scala 39:27]
  wire  _T_390; // @[LZD.scala 39:25]
  wire [1:0] _T_391; // @[Cat.scala 29:58]
  wire  _T_392; // @[Shift.scala 12:21]
  wire  _T_393; // @[Shift.scala 12:21]
  wire  _T_394; // @[LZD.scala 49:16]
  wire  _T_395; // @[LZD.scala 49:27]
  wire  _T_396; // @[LZD.scala 49:25]
  wire  _T_397; // @[LZD.scala 49:47]
  wire  _T_398; // @[LZD.scala 49:59]
  wire  _T_399; // @[LZD.scala 49:35]
  wire [2:0] _T_401; // @[Cat.scala 29:58]
  wire [3:0] _T_402; // @[LZD.scala 44:32]
  wire [1:0] _T_403; // @[LZD.scala 43:32]
  wire  _T_404; // @[LZD.scala 39:14]
  wire  _T_405; // @[LZD.scala 39:21]
  wire  _T_406; // @[LZD.scala 39:30]
  wire  _T_407; // @[LZD.scala 39:27]
  wire  _T_408; // @[LZD.scala 39:25]
  wire [1:0] _T_409; // @[Cat.scala 29:58]
  wire [1:0] _T_410; // @[LZD.scala 44:32]
  wire  _T_411; // @[LZD.scala 39:14]
  wire  _T_412; // @[LZD.scala 39:21]
  wire  _T_413; // @[LZD.scala 39:30]
  wire  _T_414; // @[LZD.scala 39:27]
  wire  _T_415; // @[LZD.scala 39:25]
  wire [1:0] _T_416; // @[Cat.scala 29:58]
  wire  _T_417; // @[Shift.scala 12:21]
  wire  _T_418; // @[Shift.scala 12:21]
  wire  _T_419; // @[LZD.scala 49:16]
  wire  _T_420; // @[LZD.scala 49:27]
  wire  _T_421; // @[LZD.scala 49:25]
  wire  _T_422; // @[LZD.scala 49:47]
  wire  _T_423; // @[LZD.scala 49:59]
  wire  _T_424; // @[LZD.scala 49:35]
  wire [2:0] _T_426; // @[Cat.scala 29:58]
  wire  _T_427; // @[Shift.scala 12:21]
  wire  _T_428; // @[Shift.scala 12:21]
  wire  _T_429; // @[LZD.scala 49:16]
  wire  _T_430; // @[LZD.scala 49:27]
  wire  _T_431; // @[LZD.scala 49:25]
  wire [1:0] _T_432; // @[LZD.scala 49:47]
  wire [1:0] _T_433; // @[LZD.scala 49:59]
  wire [1:0] _T_434; // @[LZD.scala 49:35]
  wire [3:0] _T_436; // @[Cat.scala 29:58]
  wire  _T_437; // @[Shift.scala 12:21]
  wire  _T_438; // @[Shift.scala 12:21]
  wire  _T_439; // @[LZD.scala 49:16]
  wire  _T_440; // @[LZD.scala 49:27]
  wire  _T_441; // @[LZD.scala 49:25]
  wire [2:0] _T_442; // @[LZD.scala 49:47]
  wire [2:0] _T_443; // @[LZD.scala 49:59]
  wire [2:0] _T_444; // @[LZD.scala 49:35]
  wire [4:0] _T_446; // @[Cat.scala 29:58]
  wire [13:0] _T_447; // @[LZD.scala 44:32]
  wire [7:0] _T_448; // @[LZD.scala 43:32]
  wire [3:0] _T_449; // @[LZD.scala 43:32]
  wire [1:0] _T_450; // @[LZD.scala 43:32]
  wire  _T_451; // @[LZD.scala 39:14]
  wire  _T_452; // @[LZD.scala 39:21]
  wire  _T_453; // @[LZD.scala 39:30]
  wire  _T_454; // @[LZD.scala 39:27]
  wire  _T_455; // @[LZD.scala 39:25]
  wire [1:0] _T_456; // @[Cat.scala 29:58]
  wire [1:0] _T_457; // @[LZD.scala 44:32]
  wire  _T_458; // @[LZD.scala 39:14]
  wire  _T_459; // @[LZD.scala 39:21]
  wire  _T_460; // @[LZD.scala 39:30]
  wire  _T_461; // @[LZD.scala 39:27]
  wire  _T_462; // @[LZD.scala 39:25]
  wire [1:0] _T_463; // @[Cat.scala 29:58]
  wire  _T_464; // @[Shift.scala 12:21]
  wire  _T_465; // @[Shift.scala 12:21]
  wire  _T_466; // @[LZD.scala 49:16]
  wire  _T_467; // @[LZD.scala 49:27]
  wire  _T_468; // @[LZD.scala 49:25]
  wire  _T_469; // @[LZD.scala 49:47]
  wire  _T_470; // @[LZD.scala 49:59]
  wire  _T_471; // @[LZD.scala 49:35]
  wire [2:0] _T_473; // @[Cat.scala 29:58]
  wire [3:0] _T_474; // @[LZD.scala 44:32]
  wire [1:0] _T_475; // @[LZD.scala 43:32]
  wire  _T_476; // @[LZD.scala 39:14]
  wire  _T_477; // @[LZD.scala 39:21]
  wire  _T_478; // @[LZD.scala 39:30]
  wire  _T_479; // @[LZD.scala 39:27]
  wire  _T_480; // @[LZD.scala 39:25]
  wire [1:0] _T_481; // @[Cat.scala 29:58]
  wire [1:0] _T_482; // @[LZD.scala 44:32]
  wire  _T_483; // @[LZD.scala 39:14]
  wire  _T_484; // @[LZD.scala 39:21]
  wire  _T_485; // @[LZD.scala 39:30]
  wire  _T_486; // @[LZD.scala 39:27]
  wire  _T_487; // @[LZD.scala 39:25]
  wire [1:0] _T_488; // @[Cat.scala 29:58]
  wire  _T_489; // @[Shift.scala 12:21]
  wire  _T_490; // @[Shift.scala 12:21]
  wire  _T_491; // @[LZD.scala 49:16]
  wire  _T_492; // @[LZD.scala 49:27]
  wire  _T_493; // @[LZD.scala 49:25]
  wire  _T_494; // @[LZD.scala 49:47]
  wire  _T_495; // @[LZD.scala 49:59]
  wire  _T_496; // @[LZD.scala 49:35]
  wire [2:0] _T_498; // @[Cat.scala 29:58]
  wire  _T_499; // @[Shift.scala 12:21]
  wire  _T_500; // @[Shift.scala 12:21]
  wire  _T_501; // @[LZD.scala 49:16]
  wire  _T_502; // @[LZD.scala 49:27]
  wire  _T_503; // @[LZD.scala 49:25]
  wire [1:0] _T_504; // @[LZD.scala 49:47]
  wire [1:0] _T_505; // @[LZD.scala 49:59]
  wire [1:0] _T_506; // @[LZD.scala 49:35]
  wire [3:0] _T_508; // @[Cat.scala 29:58]
  wire [5:0] _T_509; // @[LZD.scala 44:32]
  wire [3:0] _T_510; // @[LZD.scala 43:32]
  wire [1:0] _T_511; // @[LZD.scala 43:32]
  wire  _T_512; // @[LZD.scala 39:14]
  wire  _T_513; // @[LZD.scala 39:21]
  wire  _T_514; // @[LZD.scala 39:30]
  wire  _T_515; // @[LZD.scala 39:27]
  wire  _T_516; // @[LZD.scala 39:25]
  wire [1:0] _T_517; // @[Cat.scala 29:58]
  wire [1:0] _T_518; // @[LZD.scala 44:32]
  wire  _T_519; // @[LZD.scala 39:14]
  wire  _T_520; // @[LZD.scala 39:21]
  wire  _T_521; // @[LZD.scala 39:30]
  wire  _T_522; // @[LZD.scala 39:27]
  wire  _T_523; // @[LZD.scala 39:25]
  wire [1:0] _T_524; // @[Cat.scala 29:58]
  wire  _T_525; // @[Shift.scala 12:21]
  wire  _T_526; // @[Shift.scala 12:21]
  wire  _T_527; // @[LZD.scala 49:16]
  wire  _T_528; // @[LZD.scala 49:27]
  wire  _T_529; // @[LZD.scala 49:25]
  wire  _T_530; // @[LZD.scala 49:47]
  wire  _T_531; // @[LZD.scala 49:59]
  wire  _T_532; // @[LZD.scala 49:35]
  wire [2:0] _T_534; // @[Cat.scala 29:58]
  wire [1:0] _T_535; // @[LZD.scala 44:32]
  wire  _T_536; // @[LZD.scala 39:14]
  wire  _T_537; // @[LZD.scala 39:21]
  wire  _T_538; // @[LZD.scala 39:30]
  wire  _T_539; // @[LZD.scala 39:27]
  wire  _T_540; // @[LZD.scala 39:25]
  wire [1:0] _T_541; // @[Cat.scala 29:58]
  wire  _T_542; // @[Shift.scala 12:21]
  wire [1:0] _T_544; // @[LZD.scala 55:32]
  wire [1:0] _T_545; // @[LZD.scala 55:20]
  wire [2:0] _T_546; // @[Cat.scala 29:58]
  wire  _T_547; // @[Shift.scala 12:21]
  wire [2:0] _T_549; // @[LZD.scala 55:32]
  wire [2:0] _T_550; // @[LZD.scala 55:20]
  wire [3:0] _T_551; // @[Cat.scala 29:58]
  wire  _T_552; // @[Shift.scala 12:21]
  wire [3:0] _T_554; // @[LZD.scala 55:32]
  wire [3:0] _T_555; // @[LZD.scala 55:20]
  wire [4:0] _T_556; // @[Cat.scala 29:58]
  wire [4:0] _T_557; // @[convert.scala 21:22]
  wire [28:0] _T_558; // @[convert.scala 22:36]
  wire  _T_559; // @[Shift.scala 16:24]
  wire  _T_561; // @[Shift.scala 12:21]
  wire [12:0] _T_562; // @[Shift.scala 64:52]
  wire [28:0] _T_564; // @[Cat.scala 29:58]
  wire [28:0] _T_565; // @[Shift.scala 64:27]
  wire [3:0] _T_566; // @[Shift.scala 66:70]
  wire  _T_567; // @[Shift.scala 12:21]
  wire [20:0] _T_568; // @[Shift.scala 64:52]
  wire [28:0] _T_570; // @[Cat.scala 29:58]
  wire [28:0] _T_571; // @[Shift.scala 64:27]
  wire [2:0] _T_572; // @[Shift.scala 66:70]
  wire  _T_573; // @[Shift.scala 12:21]
  wire [24:0] _T_574; // @[Shift.scala 64:52]
  wire [28:0] _T_576; // @[Cat.scala 29:58]
  wire [28:0] _T_577; // @[Shift.scala 64:27]
  wire [1:0] _T_578; // @[Shift.scala 66:70]
  wire  _T_579; // @[Shift.scala 12:21]
  wire [26:0] _T_580; // @[Shift.scala 64:52]
  wire [28:0] _T_582; // @[Cat.scala 29:58]
  wire [28:0] _T_583; // @[Shift.scala 64:27]
  wire  _T_584; // @[Shift.scala 66:70]
  wire [27:0] _T_586; // @[Shift.scala 64:52]
  wire [28:0] _T_587; // @[Cat.scala 29:58]
  wire [28:0] _T_588; // @[Shift.scala 64:27]
  wire [28:0] _T_589; // @[Shift.scala 16:10]
  wire  _T_590; // @[convert.scala 23:34]
  wire [27:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_592; // @[convert.scala 25:26]
  wire [4:0] _T_594; // @[convert.scala 25:42]
  wire  _T_597; // @[convert.scala 26:67]
  wire  _T_598; // @[convert.scala 26:51]
  wire [6:0] _T_599; // @[Cat.scala 29:58]
  wire [30:0] _T_601; // @[convert.scala 29:56]
  wire  _T_602; // @[convert.scala 29:60]
  wire  _T_603; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_606; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [6:0] decB_scale; // @[convert.scala 32:24]
  wire [2:0] _T_615; // @[Bitwise.scala 71:12]
  wire  _T_616; // @[PositDivisionSqrt.scala 80:40]
  wire [34:0] sigA_S; // @[Cat.scala 29:58]
  wire  _T_619; // @[PositDivisionSqrt.scala 82:31]
  wire [34:0] sigB_S; // @[Cat.scala 29:58]
  wire  _T_622; // @[PositDivisionSqrt.scala 85:25]
  wire  invalidSqrt; // @[PositDivisionSqrt.scala 85:37]
  wire  _T_623; // @[PositDivisionSqrt.scala 88:42]
  wire  _T_624; // @[PositDivisionSqrt.scala 89:42]
  wire  _T_625; // @[PositDivisionSqrt.scala 89:56]
  wire  _T_626; // @[PositDivisionSqrt.scala 94:46]
  wire  _T_627; // @[PositDivisionSqrt.scala 94:43]
  wire  _T_628; // @[PositDivisionSqrt.scala 94:62]
  wire  _T_629; // @[PositDivisionSqrt.scala 94:59]
  wire  specialCaseA_S; // @[PositDivisionSqrt.scala 97:38]
  wire  specialCaseB_S; // @[PositDivisionSqrt.scala 98:38]
  wire  _T_630; // @[PositDivisionSqrt.scala 99:27]
  wire  _T_631; // @[PositDivisionSqrt.scala 99:46]
  wire  normalCase_S_div; // @[PositDivisionSqrt.scala 99:43]
  wire  normalCase_S_sqrt; // @[PositDivisionSqrt.scala 100:43]
  wire  normalCase_S; // @[PositDivisionSqrt.scala 101:30]
  wire [7:0] sExpQuot_S_div; // @[PositDivisionSqrt.scala 103:38]
  wire  _T_634; // @[PositDivisionSqrt.scala 104:50]
  wire  oddSqrt_S; // @[PositDivisionSqrt.scala 104:37]
  wire  idle; // @[PositDivisionSqrt.scala 109:39]
  wire  ready; // @[PositDivisionSqrt.scala 110:39]
  wire  entering; // @[PositDivisionSqrt.scala 111:35]
  wire  entering_normalCase; // @[PositDivisionSqrt.scala 112:38]
  wire  _T_635; // @[PositDivisionSqrt.scala 113:35]
  wire  _T_636; // @[PositDivisionSqrt.scala 113:58]
  wire  scaleNotChange; // @[PositDivisionSqrt.scala 113:50]
  wire  _T_637; // @[PositDivisionSqrt.scala 114:39]
  wire  skipCycle2; // @[PositDivisionSqrt.scala 114:48]
  wire  _T_638; // @[PositDivisionSqrt.scala 116:8]
  wire  _T_639; // @[PositDivisionSqrt.scala 116:14]
  wire  _T_640; // @[PositDivisionSqrt.scala 117:32]
  wire  _T_641; // @[PositDivisionSqrt.scala 117:30]
  wire [5:0] _T_643; // @[PositDivisionSqrt.scala 119:26]
  wire [5:0] _T_644; // @[PositDivisionSqrt.scala 118:20]
  wire [5:0] _GEN_9; // @[PositDivisionSqrt.scala 117:64]
  wire [5:0] _T_645; // @[PositDivisionSqrt.scala 117:64]
  wire  _T_647; // @[PositDivisionSqrt.scala 123:30]
  wire  _T_648; // @[PositDivisionSqrt.scala 123:27]
  wire [5:0] _T_650; // @[PositDivisionSqrt.scala 123:52]
  wire [5:0] _T_651; // @[PositDivisionSqrt.scala 123:20]
  wire [5:0] _T_652; // @[PositDivisionSqrt.scala 122:64]
  wire  _T_654; // @[PositDivisionSqrt.scala 124:27]
  wire [5:0] _GEN_10; // @[PositDivisionSqrt.scala 123:64]
  wire [5:0] _T_656; // @[PositDivisionSqrt.scala 123:64]
  wire [5:0] _T_657; // @[PositDivisionSqrt.scala 134:42]
  wire  _T_659; // @[PositDivisionSqrt.scala 137:31]
  wire  _T_660; // @[PositDivisionSqrt.scala 137:28]
  wire [63:0] _T_661; // @[PositDivisionSqrt.scala 146:22]
  wire [61:0] _T_662; // @[PositDivisionSqrt.scala 146:35]
  wire  _T_663; // @[PositDivisionSqrt.scala 148:26]
  wire  _T_664; // @[PositDivisionSqrt.scala 148:23]
  wire [34:0] _T_665; // @[PositDivisionSqrt.scala 148:16]
  wire  _T_666; // @[PositDivisionSqrt.scala 149:23]
  wire [35:0] _T_667; // @[PositDivisionSqrt.scala 149:46]
  wire [34:0] _T_668; // @[PositDivisionSqrt.scala 149:56]
  wire [34:0] _T_669; // @[PositDivisionSqrt.scala 149:16]
  wire [34:0] _T_670; // @[PositDivisionSqrt.scala 148:66]
  wire  _T_671; // @[PositDivisionSqrt.scala 150:17]
  wire [34:0] _T_672; // @[PositDivisionSqrt.scala 150:16]
  wire [34:0] rem; // @[PositDivisionSqrt.scala 149:66]
  wire  _T_674; // @[PositDivisionSqrt.scala 152:29]
  wire [34:0] _T_675; // @[PositDivisionSqrt.scala 152:22]
  wire  _T_676; // @[PositDivisionSqrt.scala 153:29]
  wire [31:0] _T_677; // @[PositDivisionSqrt.scala 153:22]
  wire [34:0] _GEN_11; // @[PositDivisionSqrt.scala 152:93]
  wire [34:0] _T_678; // @[PositDivisionSqrt.scala 152:93]
  wire  _T_680; // @[PositDivisionSqrt.scala 154:33]
  wire  _T_681; // @[PositDivisionSqrt.scala 154:30]
  wire  _T_682; // @[PositDivisionSqrt.scala 154:57]
  wire [34:0] _T_685; // @[Cat.scala 29:58]
  wire [34:0] _T_686; // @[PositDivisionSqrt.scala 154:22]
  wire [34:0] _T_687; // @[PositDivisionSqrt.scala 153:93]
  wire  _T_689; // @[PositDivisionSqrt.scala 155:30]
  wire  _T_690; // @[PositDivisionSqrt.scala 156:83]
  wire [30:0] _T_692; // @[Bitwise.scala 71:12]
  wire [33:0] bitMask; // @[PositDivisionSqrt.scala 145:21 PositDivisionSqrt.scala 146:14]
  wire [33:0] _GEN_12; // @[PositDivisionSqrt.scala 156:53]
  wire [33:0] _T_693; // @[PositDivisionSqrt.scala 156:53]
  wire [34:0] _GEN_13; // @[PositDivisionSqrt.scala 155:51]
  wire [34:0] _T_694; // @[PositDivisionSqrt.scala 155:51]
  wire [32:0] _T_695; // @[PositDivisionSqrt.scala 157:53]
  wire [34:0] _GEN_14; // @[PositDivisionSqrt.scala 156:89]
  wire [34:0] _T_696; // @[PositDivisionSqrt.scala 156:89]
  wire [34:0] _T_697; // @[PositDivisionSqrt.scala 155:22]
  wire [34:0] trialTerm; // @[PositDivisionSqrt.scala 154:93]
  wire  _T_699; // @[PositDivisionSqrt.scala 162:56]
  wire  _T_700; // @[PositDivisionSqrt.scala 162:40]
  wire [34:0] _T_703; // @[PositDivisionSqrt.scala 163:97]
  wire [34:0] _T_705; // @[PositDivisionSqrt.scala 164:97]
  wire [34:0] _T_706; // @[PositDivisionSqrt.scala 161:92]
  wire [35:0] _T_711; // @[PositDivisionSqrt.scala 168:98]
  wire [34:0] _T_712; // @[PositDivisionSqrt.scala 168:108]
  wire [34:0] _T_714; // @[PositDivisionSqrt.scala 168:112]
  wire [34:0] _T_718; // @[PositDivisionSqrt.scala 169:112]
  wire [34:0] _T_719; // @[PositDivisionSqrt.scala 166:26]
  wire [34:0] trialRem; // @[PositDivisionSqrt.scala 159:27]
  wire  _T_720; // @[PositDivisionSqrt.scala 173:35]
  wire  trIsZero; // @[PositDivisionSqrt.scala 173:25]
  wire  _T_721; // @[PositDivisionSqrt.scala 174:30]
  wire  remIsZero; // @[PositDivisionSqrt.scala 174:25]
  wire  _T_723; // @[PositDivisionSqrt.scala 176:64]
  wire  _T_724; // @[PositDivisionSqrt.scala 176:49]
  wire  _T_725; // @[PositDivisionSqrt.scala 176:29]
  wire  _T_726; // @[PositDivisionSqrt.scala 178:61]
  wire  _T_727; // @[PositDivisionSqrt.scala 178:49]
  wire  _T_729; // @[Mux.scala 87:16]
  wire  newBit; // @[Mux.scala 87:16]
  wire  _T_730; // @[PositDivisionSqrt.scala 183:41]
  wire  _T_731; // @[PositDivisionSqrt.scala 183:51]
  wire  _T_732; // @[PositDivisionSqrt.scala 183:48]
  wire  _T_733; // @[PositDivisionSqrt.scala 183:28]
  wire  _T_736; // @[PositDivisionSqrt.scala 187:39]
  wire  _T_737; // @[PositDivisionSqrt.scala 187:28]
  wire [34:0] _T_740; // @[PositDivisionSqrt.scala 188:47]
  wire [34:0] _T_741; // @[PositDivisionSqrt.scala 188:18]
  wire [32:0] _T_743; // @[PositDivisionSqrt.scala 189:18]
  wire [34:0] _GEN_15; // @[PositDivisionSqrt.scala 188:78]
  wire [34:0] _T_744; // @[PositDivisionSqrt.scala 188:78]
  wire [34:0] _GEN_16; // @[PositDivisionSqrt.scala 190:47]
  wire [34:0] _T_746; // @[PositDivisionSqrt.scala 190:47]
  wire [34:0] _T_747; // @[PositDivisionSqrt.scala 190:18]
  wire [34:0] _T_748; // @[PositDivisionSqrt.scala 189:78]
  wire [1:0] _T_750; // @[PositDivisionSqrt.scala 196:53]
  wire [1:0] sigXBias; // @[PositDivisionSqrt.scala 196:21]
  wire [34:0] _GEN_17; // @[PositDivisionSqrt.scala 197:25]
  wire [34:0] realSigX; // @[PositDivisionSqrt.scala 197:25]
  wire [27:0] _T_753; // @[PositDivisionSqrt.scala 200:97]
  wire [27:0] _T_754; // @[PositDivisionSqrt.scala 201:97]
  wire [27:0] realFrac; // @[PositDivisionSqrt.scala 198:21]
  wire  _T_755; // @[PositDivisionSqrt.scala 205:33]
  wire  _T_756; // @[PositDivisionSqrt.scala 205:58]
  wire  _T_757; // @[PositDivisionSqrt.scala 205:48]
  wire  scaleNeedSub; // @[PositDivisionSqrt.scala 205:23]
  wire  _T_759; // @[PositDivisionSqrt.scala 206:56]
  wire  notNeedSubTwo; // @[PositDivisionSqrt.scala 206:46]
  wire  scaleSubOne; // @[PositDivisionSqrt.scala 207:36]
  wire  _T_760; // @[PositDivisionSqrt.scala 208:38]
  wire  scaleSubTwo; // @[PositDivisionSqrt.scala 208:36]
  wire [1:0] _T_761; // @[Cat.scala 29:58]
  wire [2:0] _T_762; // @[PositDivisionSqrt.scala 209:63]
  wire [7:0] _GEN_18; // @[PositDivisionSqrt.scala 209:31]
  wire [7:0] _T_764; // @[PositDivisionSqrt.scala 209:31]
  wire [7:0] realExp; // @[PositDivisionSqrt.scala 209:31]
  wire  underflow; // @[PositDivisionSqrt.scala 210:31]
  wire  overflow; // @[PositDivisionSqrt.scala 211:31]
  wire  decQ_sign; // @[PositDivisionSqrt.scala 215:33]
  wire [7:0] _T_766; // @[Mux.scala 87:16]
  wire [7:0] _T_767; // @[Mux.scala 87:16]
  wire [2:0] _T_768; // @[PositDivisionSqrt.scala 224:48]
  wire [2:0] _T_769; // @[PositDivisionSqrt.scala 224:64]
  wire [2:0] decQ_grs; // @[PositDivisionSqrt.scala 224:23]
  wire  outValid; // @[PositDivisionSqrt.scala 229:28]
  wire [6:0] _GEN_19; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire [6:0] decQ_scale; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire  _T_775; // @[convert.scala 46:61]
  wire  _T_776; // @[convert.scala 46:52]
  wire  _T_778; // @[convert.scala 46:42]
  wire [5:0] _T_779; // @[convert.scala 48:34]
  wire  _T_780; // @[convert.scala 49:36]
  wire [5:0] _T_782; // @[convert.scala 50:36]
  wire [5:0] _T_783; // @[convert.scala 50:36]
  wire [5:0] _T_784; // @[convert.scala 50:28]
  wire  _T_785; // @[convert.scala 51:31]
  wire  _T_786; // @[convert.scala 52:43]
  wire [33:0] _T_790; // @[Cat.scala 29:58]
  wire [5:0] _T_791; // @[Shift.scala 39:17]
  wire  _T_792; // @[Shift.scala 39:24]
  wire [1:0] _T_794; // @[Shift.scala 90:30]
  wire [31:0] _T_795; // @[Shift.scala 90:48]
  wire  _T_796; // @[Shift.scala 90:57]
  wire [1:0] _GEN_20; // @[Shift.scala 90:39]
  wire [1:0] _T_797; // @[Shift.scala 90:39]
  wire  _T_798; // @[Shift.scala 12:21]
  wire  _T_799; // @[Shift.scala 12:21]
  wire [31:0] _T_801; // @[Bitwise.scala 71:12]
  wire [33:0] _T_802; // @[Cat.scala 29:58]
  wire [33:0] _T_803; // @[Shift.scala 91:22]
  wire [4:0] _T_804; // @[Shift.scala 92:77]
  wire [17:0] _T_805; // @[Shift.scala 90:30]
  wire [15:0] _T_806; // @[Shift.scala 90:48]
  wire  _T_807; // @[Shift.scala 90:57]
  wire [17:0] _GEN_21; // @[Shift.scala 90:39]
  wire [17:0] _T_808; // @[Shift.scala 90:39]
  wire  _T_809; // @[Shift.scala 12:21]
  wire  _T_810; // @[Shift.scala 12:21]
  wire [15:0] _T_812; // @[Bitwise.scala 71:12]
  wire [33:0] _T_813; // @[Cat.scala 29:58]
  wire [33:0] _T_814; // @[Shift.scala 91:22]
  wire [3:0] _T_815; // @[Shift.scala 92:77]
  wire [25:0] _T_816; // @[Shift.scala 90:30]
  wire [7:0] _T_817; // @[Shift.scala 90:48]
  wire  _T_818; // @[Shift.scala 90:57]
  wire [25:0] _GEN_22; // @[Shift.scala 90:39]
  wire [25:0] _T_819; // @[Shift.scala 90:39]
  wire  _T_820; // @[Shift.scala 12:21]
  wire  _T_821; // @[Shift.scala 12:21]
  wire [7:0] _T_823; // @[Bitwise.scala 71:12]
  wire [33:0] _T_824; // @[Cat.scala 29:58]
  wire [33:0] _T_825; // @[Shift.scala 91:22]
  wire [2:0] _T_826; // @[Shift.scala 92:77]
  wire [29:0] _T_827; // @[Shift.scala 90:30]
  wire [3:0] _T_828; // @[Shift.scala 90:48]
  wire  _T_829; // @[Shift.scala 90:57]
  wire [29:0] _GEN_23; // @[Shift.scala 90:39]
  wire [29:0] _T_830; // @[Shift.scala 90:39]
  wire  _T_831; // @[Shift.scala 12:21]
  wire  _T_832; // @[Shift.scala 12:21]
  wire [3:0] _T_834; // @[Bitwise.scala 71:12]
  wire [33:0] _T_835; // @[Cat.scala 29:58]
  wire [33:0] _T_836; // @[Shift.scala 91:22]
  wire [1:0] _T_837; // @[Shift.scala 92:77]
  wire [31:0] _T_838; // @[Shift.scala 90:30]
  wire [1:0] _T_839; // @[Shift.scala 90:48]
  wire  _T_840; // @[Shift.scala 90:57]
  wire [31:0] _GEN_24; // @[Shift.scala 90:39]
  wire [31:0] _T_841; // @[Shift.scala 90:39]
  wire  _T_842; // @[Shift.scala 12:21]
  wire  _T_843; // @[Shift.scala 12:21]
  wire [1:0] _T_845; // @[Bitwise.scala 71:12]
  wire [33:0] _T_846; // @[Cat.scala 29:58]
  wire [33:0] _T_847; // @[Shift.scala 91:22]
  wire  _T_848; // @[Shift.scala 92:77]
  wire [32:0] _T_849; // @[Shift.scala 90:30]
  wire  _T_850; // @[Shift.scala 90:48]
  wire [32:0] _GEN_25; // @[Shift.scala 90:39]
  wire [32:0] _T_852; // @[Shift.scala 90:39]
  wire  _T_854; // @[Shift.scala 12:21]
  wire [33:0] _T_855; // @[Cat.scala 29:58]
  wire [33:0] _T_856; // @[Shift.scala 91:22]
  wire [33:0] _T_859; // @[Bitwise.scala 71:12]
  wire [33:0] _T_860; // @[Shift.scala 39:10]
  wire  _T_861; // @[convert.scala 55:31]
  wire  _T_862; // @[convert.scala 56:31]
  wire  _T_863; // @[convert.scala 57:31]
  wire  _T_864; // @[convert.scala 58:31]
  wire [30:0] _T_865; // @[convert.scala 59:69]
  wire  _T_866; // @[convert.scala 59:81]
  wire  _T_867; // @[convert.scala 59:50]
  wire  _T_869; // @[convert.scala 60:81]
  wire  _T_870; // @[convert.scala 61:44]
  wire  _T_871; // @[convert.scala 61:52]
  wire  _T_872; // @[convert.scala 61:36]
  wire  _T_873; // @[convert.scala 62:63]
  wire  _T_874; // @[convert.scala 62:103]
  wire  _T_875; // @[convert.scala 62:60]
  wire [30:0] _GEN_26; // @[convert.scala 63:56]
  wire [30:0] _T_878; // @[convert.scala 63:56]
  wire [31:0] _T_879; // @[Cat.scala 29:58]
  wire [31:0] _T_881; // @[Mux.scala 87:16]
  assign _T_1 = io_A[31]; // @[convert.scala 18:24]
  assign _T_2 = io_A[30]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[30:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[29:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[29:14]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[15:8]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8[7:4]; // @[LZD.scala 43:32]
  assign _T_10 = _T_9[3:2]; // @[LZD.scala 43:32]
  assign _T_11 = _T_10 != 2'h0; // @[LZD.scala 39:14]
  assign _T_12 = _T_10[1]; // @[LZD.scala 39:21]
  assign _T_13 = _T_10[0]; // @[LZD.scala 39:30]
  assign _T_14 = ~ _T_13; // @[LZD.scala 39:27]
  assign _T_15 = _T_12 | _T_14; // @[LZD.scala 39:25]
  assign _T_16 = {_T_11,_T_15}; // @[Cat.scala 29:58]
  assign _T_17 = _T_9[1:0]; // @[LZD.scala 44:32]
  assign _T_18 = _T_17 != 2'h0; // @[LZD.scala 39:14]
  assign _T_19 = _T_17[1]; // @[LZD.scala 39:21]
  assign _T_20 = _T_17[0]; // @[LZD.scala 39:30]
  assign _T_21 = ~ _T_20; // @[LZD.scala 39:27]
  assign _T_22 = _T_19 | _T_21; // @[LZD.scala 39:25]
  assign _T_23 = {_T_18,_T_22}; // @[Cat.scala 29:58]
  assign _T_24 = _T_16[1]; // @[Shift.scala 12:21]
  assign _T_25 = _T_23[1]; // @[Shift.scala 12:21]
  assign _T_26 = _T_24 | _T_25; // @[LZD.scala 49:16]
  assign _T_27 = ~ _T_25; // @[LZD.scala 49:27]
  assign _T_28 = _T_24 | _T_27; // @[LZD.scala 49:25]
  assign _T_29 = _T_16[0:0]; // @[LZD.scala 49:47]
  assign _T_30 = _T_23[0:0]; // @[LZD.scala 49:59]
  assign _T_31 = _T_24 ? _T_29 : _T_30; // @[LZD.scala 49:35]
  assign _T_33 = {_T_26,_T_28,_T_31}; // @[Cat.scala 29:58]
  assign _T_34 = _T_8[3:0]; // @[LZD.scala 44:32]
  assign _T_35 = _T_34[3:2]; // @[LZD.scala 43:32]
  assign _T_36 = _T_35 != 2'h0; // @[LZD.scala 39:14]
  assign _T_37 = _T_35[1]; // @[LZD.scala 39:21]
  assign _T_38 = _T_35[0]; // @[LZD.scala 39:30]
  assign _T_39 = ~ _T_38; // @[LZD.scala 39:27]
  assign _T_40 = _T_37 | _T_39; // @[LZD.scala 39:25]
  assign _T_41 = {_T_36,_T_40}; // @[Cat.scala 29:58]
  assign _T_42 = _T_34[1:0]; // @[LZD.scala 44:32]
  assign _T_43 = _T_42 != 2'h0; // @[LZD.scala 39:14]
  assign _T_44 = _T_42[1]; // @[LZD.scala 39:21]
  assign _T_45 = _T_42[0]; // @[LZD.scala 39:30]
  assign _T_46 = ~ _T_45; // @[LZD.scala 39:27]
  assign _T_47 = _T_44 | _T_46; // @[LZD.scala 39:25]
  assign _T_48 = {_T_43,_T_47}; // @[Cat.scala 29:58]
  assign _T_49 = _T_41[1]; // @[Shift.scala 12:21]
  assign _T_50 = _T_48[1]; // @[Shift.scala 12:21]
  assign _T_51 = _T_49 | _T_50; // @[LZD.scala 49:16]
  assign _T_52 = ~ _T_50; // @[LZD.scala 49:27]
  assign _T_53 = _T_49 | _T_52; // @[LZD.scala 49:25]
  assign _T_54 = _T_41[0:0]; // @[LZD.scala 49:47]
  assign _T_55 = _T_48[0:0]; // @[LZD.scala 49:59]
  assign _T_56 = _T_49 ? _T_54 : _T_55; // @[LZD.scala 49:35]
  assign _T_58 = {_T_51,_T_53,_T_56}; // @[Cat.scala 29:58]
  assign _T_59 = _T_33[2]; // @[Shift.scala 12:21]
  assign _T_60 = _T_58[2]; // @[Shift.scala 12:21]
  assign _T_61 = _T_59 | _T_60; // @[LZD.scala 49:16]
  assign _T_62 = ~ _T_60; // @[LZD.scala 49:27]
  assign _T_63 = _T_59 | _T_62; // @[LZD.scala 49:25]
  assign _T_64 = _T_33[1:0]; // @[LZD.scala 49:47]
  assign _T_65 = _T_58[1:0]; // @[LZD.scala 49:59]
  assign _T_66 = _T_59 ? _T_64 : _T_65; // @[LZD.scala 49:35]
  assign _T_68 = {_T_61,_T_63,_T_66}; // @[Cat.scala 29:58]
  assign _T_69 = _T_7[7:0]; // @[LZD.scala 44:32]
  assign _T_70 = _T_69[7:4]; // @[LZD.scala 43:32]
  assign _T_71 = _T_70[3:2]; // @[LZD.scala 43:32]
  assign _T_72 = _T_71 != 2'h0; // @[LZD.scala 39:14]
  assign _T_73 = _T_71[1]; // @[LZD.scala 39:21]
  assign _T_74 = _T_71[0]; // @[LZD.scala 39:30]
  assign _T_75 = ~ _T_74; // @[LZD.scala 39:27]
  assign _T_76 = _T_73 | _T_75; // @[LZD.scala 39:25]
  assign _T_77 = {_T_72,_T_76}; // @[Cat.scala 29:58]
  assign _T_78 = _T_70[1:0]; // @[LZD.scala 44:32]
  assign _T_79 = _T_78 != 2'h0; // @[LZD.scala 39:14]
  assign _T_80 = _T_78[1]; // @[LZD.scala 39:21]
  assign _T_81 = _T_78[0]; // @[LZD.scala 39:30]
  assign _T_82 = ~ _T_81; // @[LZD.scala 39:27]
  assign _T_83 = _T_80 | _T_82; // @[LZD.scala 39:25]
  assign _T_84 = {_T_79,_T_83}; // @[Cat.scala 29:58]
  assign _T_85 = _T_77[1]; // @[Shift.scala 12:21]
  assign _T_86 = _T_84[1]; // @[Shift.scala 12:21]
  assign _T_87 = _T_85 | _T_86; // @[LZD.scala 49:16]
  assign _T_88 = ~ _T_86; // @[LZD.scala 49:27]
  assign _T_89 = _T_85 | _T_88; // @[LZD.scala 49:25]
  assign _T_90 = _T_77[0:0]; // @[LZD.scala 49:47]
  assign _T_91 = _T_84[0:0]; // @[LZD.scala 49:59]
  assign _T_92 = _T_85 ? _T_90 : _T_91; // @[LZD.scala 49:35]
  assign _T_94 = {_T_87,_T_89,_T_92}; // @[Cat.scala 29:58]
  assign _T_95 = _T_69[3:0]; // @[LZD.scala 44:32]
  assign _T_96 = _T_95[3:2]; // @[LZD.scala 43:32]
  assign _T_97 = _T_96 != 2'h0; // @[LZD.scala 39:14]
  assign _T_98 = _T_96[1]; // @[LZD.scala 39:21]
  assign _T_99 = _T_96[0]; // @[LZD.scala 39:30]
  assign _T_100 = ~ _T_99; // @[LZD.scala 39:27]
  assign _T_101 = _T_98 | _T_100; // @[LZD.scala 39:25]
  assign _T_102 = {_T_97,_T_101}; // @[Cat.scala 29:58]
  assign _T_103 = _T_95[1:0]; // @[LZD.scala 44:32]
  assign _T_104 = _T_103 != 2'h0; // @[LZD.scala 39:14]
  assign _T_105 = _T_103[1]; // @[LZD.scala 39:21]
  assign _T_106 = _T_103[0]; // @[LZD.scala 39:30]
  assign _T_107 = ~ _T_106; // @[LZD.scala 39:27]
  assign _T_108 = _T_105 | _T_107; // @[LZD.scala 39:25]
  assign _T_109 = {_T_104,_T_108}; // @[Cat.scala 29:58]
  assign _T_110 = _T_102[1]; // @[Shift.scala 12:21]
  assign _T_111 = _T_109[1]; // @[Shift.scala 12:21]
  assign _T_112 = _T_110 | _T_111; // @[LZD.scala 49:16]
  assign _T_113 = ~ _T_111; // @[LZD.scala 49:27]
  assign _T_114 = _T_110 | _T_113; // @[LZD.scala 49:25]
  assign _T_115 = _T_102[0:0]; // @[LZD.scala 49:47]
  assign _T_116 = _T_109[0:0]; // @[LZD.scala 49:59]
  assign _T_117 = _T_110 ? _T_115 : _T_116; // @[LZD.scala 49:35]
  assign _T_119 = {_T_112,_T_114,_T_117}; // @[Cat.scala 29:58]
  assign _T_120 = _T_94[2]; // @[Shift.scala 12:21]
  assign _T_121 = _T_119[2]; // @[Shift.scala 12:21]
  assign _T_122 = _T_120 | _T_121; // @[LZD.scala 49:16]
  assign _T_123 = ~ _T_121; // @[LZD.scala 49:27]
  assign _T_124 = _T_120 | _T_123; // @[LZD.scala 49:25]
  assign _T_125 = _T_94[1:0]; // @[LZD.scala 49:47]
  assign _T_126 = _T_119[1:0]; // @[LZD.scala 49:59]
  assign _T_127 = _T_120 ? _T_125 : _T_126; // @[LZD.scala 49:35]
  assign _T_129 = {_T_122,_T_124,_T_127}; // @[Cat.scala 29:58]
  assign _T_130 = _T_68[3]; // @[Shift.scala 12:21]
  assign _T_131 = _T_129[3]; // @[Shift.scala 12:21]
  assign _T_132 = _T_130 | _T_131; // @[LZD.scala 49:16]
  assign _T_133 = ~ _T_131; // @[LZD.scala 49:27]
  assign _T_134 = _T_130 | _T_133; // @[LZD.scala 49:25]
  assign _T_135 = _T_68[2:0]; // @[LZD.scala 49:47]
  assign _T_136 = _T_129[2:0]; // @[LZD.scala 49:59]
  assign _T_137 = _T_130 ? _T_135 : _T_136; // @[LZD.scala 49:35]
  assign _T_139 = {_T_132,_T_134,_T_137}; // @[Cat.scala 29:58]
  assign _T_140 = _T_6[13:0]; // @[LZD.scala 44:32]
  assign _T_141 = _T_140[13:6]; // @[LZD.scala 43:32]
  assign _T_142 = _T_141[7:4]; // @[LZD.scala 43:32]
  assign _T_143 = _T_142[3:2]; // @[LZD.scala 43:32]
  assign _T_144 = _T_143 != 2'h0; // @[LZD.scala 39:14]
  assign _T_145 = _T_143[1]; // @[LZD.scala 39:21]
  assign _T_146 = _T_143[0]; // @[LZD.scala 39:30]
  assign _T_147 = ~ _T_146; // @[LZD.scala 39:27]
  assign _T_148 = _T_145 | _T_147; // @[LZD.scala 39:25]
  assign _T_149 = {_T_144,_T_148}; // @[Cat.scala 29:58]
  assign _T_150 = _T_142[1:0]; // @[LZD.scala 44:32]
  assign _T_151 = _T_150 != 2'h0; // @[LZD.scala 39:14]
  assign _T_152 = _T_150[1]; // @[LZD.scala 39:21]
  assign _T_153 = _T_150[0]; // @[LZD.scala 39:30]
  assign _T_154 = ~ _T_153; // @[LZD.scala 39:27]
  assign _T_155 = _T_152 | _T_154; // @[LZD.scala 39:25]
  assign _T_156 = {_T_151,_T_155}; // @[Cat.scala 29:58]
  assign _T_157 = _T_149[1]; // @[Shift.scala 12:21]
  assign _T_158 = _T_156[1]; // @[Shift.scala 12:21]
  assign _T_159 = _T_157 | _T_158; // @[LZD.scala 49:16]
  assign _T_160 = ~ _T_158; // @[LZD.scala 49:27]
  assign _T_161 = _T_157 | _T_160; // @[LZD.scala 49:25]
  assign _T_162 = _T_149[0:0]; // @[LZD.scala 49:47]
  assign _T_163 = _T_156[0:0]; // @[LZD.scala 49:59]
  assign _T_164 = _T_157 ? _T_162 : _T_163; // @[LZD.scala 49:35]
  assign _T_166 = {_T_159,_T_161,_T_164}; // @[Cat.scala 29:58]
  assign _T_167 = _T_141[3:0]; // @[LZD.scala 44:32]
  assign _T_168 = _T_167[3:2]; // @[LZD.scala 43:32]
  assign _T_169 = _T_168 != 2'h0; // @[LZD.scala 39:14]
  assign _T_170 = _T_168[1]; // @[LZD.scala 39:21]
  assign _T_171 = _T_168[0]; // @[LZD.scala 39:30]
  assign _T_172 = ~ _T_171; // @[LZD.scala 39:27]
  assign _T_173 = _T_170 | _T_172; // @[LZD.scala 39:25]
  assign _T_174 = {_T_169,_T_173}; // @[Cat.scala 29:58]
  assign _T_175 = _T_167[1:0]; // @[LZD.scala 44:32]
  assign _T_176 = _T_175 != 2'h0; // @[LZD.scala 39:14]
  assign _T_177 = _T_175[1]; // @[LZD.scala 39:21]
  assign _T_178 = _T_175[0]; // @[LZD.scala 39:30]
  assign _T_179 = ~ _T_178; // @[LZD.scala 39:27]
  assign _T_180 = _T_177 | _T_179; // @[LZD.scala 39:25]
  assign _T_181 = {_T_176,_T_180}; // @[Cat.scala 29:58]
  assign _T_182 = _T_174[1]; // @[Shift.scala 12:21]
  assign _T_183 = _T_181[1]; // @[Shift.scala 12:21]
  assign _T_184 = _T_182 | _T_183; // @[LZD.scala 49:16]
  assign _T_185 = ~ _T_183; // @[LZD.scala 49:27]
  assign _T_186 = _T_182 | _T_185; // @[LZD.scala 49:25]
  assign _T_187 = _T_174[0:0]; // @[LZD.scala 49:47]
  assign _T_188 = _T_181[0:0]; // @[LZD.scala 49:59]
  assign _T_189 = _T_182 ? _T_187 : _T_188; // @[LZD.scala 49:35]
  assign _T_191 = {_T_184,_T_186,_T_189}; // @[Cat.scala 29:58]
  assign _T_192 = _T_166[2]; // @[Shift.scala 12:21]
  assign _T_193 = _T_191[2]; // @[Shift.scala 12:21]
  assign _T_194 = _T_192 | _T_193; // @[LZD.scala 49:16]
  assign _T_195 = ~ _T_193; // @[LZD.scala 49:27]
  assign _T_196 = _T_192 | _T_195; // @[LZD.scala 49:25]
  assign _T_197 = _T_166[1:0]; // @[LZD.scala 49:47]
  assign _T_198 = _T_191[1:0]; // @[LZD.scala 49:59]
  assign _T_199 = _T_192 ? _T_197 : _T_198; // @[LZD.scala 49:35]
  assign _T_201 = {_T_194,_T_196,_T_199}; // @[Cat.scala 29:58]
  assign _T_202 = _T_140[5:0]; // @[LZD.scala 44:32]
  assign _T_203 = _T_202[5:2]; // @[LZD.scala 43:32]
  assign _T_204 = _T_203[3:2]; // @[LZD.scala 43:32]
  assign _T_205 = _T_204 != 2'h0; // @[LZD.scala 39:14]
  assign _T_206 = _T_204[1]; // @[LZD.scala 39:21]
  assign _T_207 = _T_204[0]; // @[LZD.scala 39:30]
  assign _T_208 = ~ _T_207; // @[LZD.scala 39:27]
  assign _T_209 = _T_206 | _T_208; // @[LZD.scala 39:25]
  assign _T_210 = {_T_205,_T_209}; // @[Cat.scala 29:58]
  assign _T_211 = _T_203[1:0]; // @[LZD.scala 44:32]
  assign _T_212 = _T_211 != 2'h0; // @[LZD.scala 39:14]
  assign _T_213 = _T_211[1]; // @[LZD.scala 39:21]
  assign _T_214 = _T_211[0]; // @[LZD.scala 39:30]
  assign _T_215 = ~ _T_214; // @[LZD.scala 39:27]
  assign _T_216 = _T_213 | _T_215; // @[LZD.scala 39:25]
  assign _T_217 = {_T_212,_T_216}; // @[Cat.scala 29:58]
  assign _T_218 = _T_210[1]; // @[Shift.scala 12:21]
  assign _T_219 = _T_217[1]; // @[Shift.scala 12:21]
  assign _T_220 = _T_218 | _T_219; // @[LZD.scala 49:16]
  assign _T_221 = ~ _T_219; // @[LZD.scala 49:27]
  assign _T_222 = _T_218 | _T_221; // @[LZD.scala 49:25]
  assign _T_223 = _T_210[0:0]; // @[LZD.scala 49:47]
  assign _T_224 = _T_217[0:0]; // @[LZD.scala 49:59]
  assign _T_225 = _T_218 ? _T_223 : _T_224; // @[LZD.scala 49:35]
  assign _T_227 = {_T_220,_T_222,_T_225}; // @[Cat.scala 29:58]
  assign _T_228 = _T_202[1:0]; // @[LZD.scala 44:32]
  assign _T_229 = _T_228 != 2'h0; // @[LZD.scala 39:14]
  assign _T_230 = _T_228[1]; // @[LZD.scala 39:21]
  assign _T_231 = _T_228[0]; // @[LZD.scala 39:30]
  assign _T_232 = ~ _T_231; // @[LZD.scala 39:27]
  assign _T_233 = _T_230 | _T_232; // @[LZD.scala 39:25]
  assign _T_234 = {_T_229,_T_233}; // @[Cat.scala 29:58]
  assign _T_235 = _T_227[2]; // @[Shift.scala 12:21]
  assign _T_237 = _T_227[1:0]; // @[LZD.scala 55:32]
  assign _T_238 = _T_235 ? _T_237 : _T_234; // @[LZD.scala 55:20]
  assign _T_239 = {_T_235,_T_238}; // @[Cat.scala 29:58]
  assign _T_240 = _T_201[3]; // @[Shift.scala 12:21]
  assign _T_242 = _T_201[2:0]; // @[LZD.scala 55:32]
  assign _T_243 = _T_240 ? _T_242 : _T_239; // @[LZD.scala 55:20]
  assign _T_244 = {_T_240,_T_243}; // @[Cat.scala 29:58]
  assign _T_245 = _T_139[4]; // @[Shift.scala 12:21]
  assign _T_247 = _T_139[3:0]; // @[LZD.scala 55:32]
  assign _T_248 = _T_245 ? _T_247 : _T_244; // @[LZD.scala 55:20]
  assign _T_249 = {_T_245,_T_248}; // @[Cat.scala 29:58]
  assign _T_250 = ~ _T_249; // @[convert.scala 21:22]
  assign _T_251 = io_A[28:0]; // @[convert.scala 22:36]
  assign _T_252 = _T_250 < 5'h1d; // @[Shift.scala 16:24]
  assign _T_254 = _T_250[4]; // @[Shift.scala 12:21]
  assign _T_255 = _T_251[12:0]; // @[Shift.scala 64:52]
  assign _T_257 = {_T_255,16'h0}; // @[Cat.scala 29:58]
  assign _T_258 = _T_254 ? _T_257 : _T_251; // @[Shift.scala 64:27]
  assign _T_259 = _T_250[3:0]; // @[Shift.scala 66:70]
  assign _T_260 = _T_259[3]; // @[Shift.scala 12:21]
  assign _T_261 = _T_258[20:0]; // @[Shift.scala 64:52]
  assign _T_263 = {_T_261,8'h0}; // @[Cat.scala 29:58]
  assign _T_264 = _T_260 ? _T_263 : _T_258; // @[Shift.scala 64:27]
  assign _T_265 = _T_259[2:0]; // @[Shift.scala 66:70]
  assign _T_266 = _T_265[2]; // @[Shift.scala 12:21]
  assign _T_267 = _T_264[24:0]; // @[Shift.scala 64:52]
  assign _T_269 = {_T_267,4'h0}; // @[Cat.scala 29:58]
  assign _T_270 = _T_266 ? _T_269 : _T_264; // @[Shift.scala 64:27]
  assign _T_271 = _T_265[1:0]; // @[Shift.scala 66:70]
  assign _T_272 = _T_271[1]; // @[Shift.scala 12:21]
  assign _T_273 = _T_270[26:0]; // @[Shift.scala 64:52]
  assign _T_275 = {_T_273,2'h0}; // @[Cat.scala 29:58]
  assign _T_276 = _T_272 ? _T_275 : _T_270; // @[Shift.scala 64:27]
  assign _T_277 = _T_271[0:0]; // @[Shift.scala 66:70]
  assign _T_279 = _T_276[27:0]; // @[Shift.scala 64:52]
  assign _T_280 = {_T_279,1'h0}; // @[Cat.scala 29:58]
  assign _T_281 = _T_277 ? _T_280 : _T_276; // @[Shift.scala 64:27]
  assign _T_282 = _T_252 ? _T_281 : 29'h0; // @[Shift.scala 16:10]
  assign _T_283 = _T_282[28:28]; // @[convert.scala 23:34]
  assign decA_fraction = _T_282[27:0]; // @[convert.scala 24:34]
  assign _T_285 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_287 = _T_3 ? _T_250 : _T_249; // @[convert.scala 25:42]
  assign _T_290 = ~ _T_283; // @[convert.scala 26:67]
  assign _T_291 = _T_1 ? _T_290 : _T_283; // @[convert.scala 26:51]
  assign _T_292 = {_T_285,_T_287,_T_291}; // @[Cat.scala 29:58]
  assign _T_294 = io_A[30:0]; // @[convert.scala 29:56]
  assign _T_295 = _T_294 != 31'h0; // @[convert.scala 29:60]
  assign _T_296 = ~ _T_295; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_296; // @[convert.scala 29:39]
  assign _T_299 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_299 & _T_296; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_292); // @[convert.scala 32:24]
  assign _T_308 = io_B[31]; // @[convert.scala 18:24]
  assign _T_309 = io_B[30]; // @[convert.scala 18:40]
  assign _T_310 = _T_308 ^ _T_309; // @[convert.scala 18:36]
  assign _T_311 = io_B[30:1]; // @[convert.scala 19:24]
  assign _T_312 = io_B[29:0]; // @[convert.scala 19:43]
  assign _T_313 = _T_311 ^ _T_312; // @[convert.scala 19:39]
  assign _T_314 = _T_313[29:14]; // @[LZD.scala 43:32]
  assign _T_315 = _T_314[15:8]; // @[LZD.scala 43:32]
  assign _T_316 = _T_315[7:4]; // @[LZD.scala 43:32]
  assign _T_317 = _T_316[3:2]; // @[LZD.scala 43:32]
  assign _T_318 = _T_317 != 2'h0; // @[LZD.scala 39:14]
  assign _T_319 = _T_317[1]; // @[LZD.scala 39:21]
  assign _T_320 = _T_317[0]; // @[LZD.scala 39:30]
  assign _T_321 = ~ _T_320; // @[LZD.scala 39:27]
  assign _T_322 = _T_319 | _T_321; // @[LZD.scala 39:25]
  assign _T_323 = {_T_318,_T_322}; // @[Cat.scala 29:58]
  assign _T_324 = _T_316[1:0]; // @[LZD.scala 44:32]
  assign _T_325 = _T_324 != 2'h0; // @[LZD.scala 39:14]
  assign _T_326 = _T_324[1]; // @[LZD.scala 39:21]
  assign _T_327 = _T_324[0]; // @[LZD.scala 39:30]
  assign _T_328 = ~ _T_327; // @[LZD.scala 39:27]
  assign _T_329 = _T_326 | _T_328; // @[LZD.scala 39:25]
  assign _T_330 = {_T_325,_T_329}; // @[Cat.scala 29:58]
  assign _T_331 = _T_323[1]; // @[Shift.scala 12:21]
  assign _T_332 = _T_330[1]; // @[Shift.scala 12:21]
  assign _T_333 = _T_331 | _T_332; // @[LZD.scala 49:16]
  assign _T_334 = ~ _T_332; // @[LZD.scala 49:27]
  assign _T_335 = _T_331 | _T_334; // @[LZD.scala 49:25]
  assign _T_336 = _T_323[0:0]; // @[LZD.scala 49:47]
  assign _T_337 = _T_330[0:0]; // @[LZD.scala 49:59]
  assign _T_338 = _T_331 ? _T_336 : _T_337; // @[LZD.scala 49:35]
  assign _T_340 = {_T_333,_T_335,_T_338}; // @[Cat.scala 29:58]
  assign _T_341 = _T_315[3:0]; // @[LZD.scala 44:32]
  assign _T_342 = _T_341[3:2]; // @[LZD.scala 43:32]
  assign _T_343 = _T_342 != 2'h0; // @[LZD.scala 39:14]
  assign _T_344 = _T_342[1]; // @[LZD.scala 39:21]
  assign _T_345 = _T_342[0]; // @[LZD.scala 39:30]
  assign _T_346 = ~ _T_345; // @[LZD.scala 39:27]
  assign _T_347 = _T_344 | _T_346; // @[LZD.scala 39:25]
  assign _T_348 = {_T_343,_T_347}; // @[Cat.scala 29:58]
  assign _T_349 = _T_341[1:0]; // @[LZD.scala 44:32]
  assign _T_350 = _T_349 != 2'h0; // @[LZD.scala 39:14]
  assign _T_351 = _T_349[1]; // @[LZD.scala 39:21]
  assign _T_352 = _T_349[0]; // @[LZD.scala 39:30]
  assign _T_353 = ~ _T_352; // @[LZD.scala 39:27]
  assign _T_354 = _T_351 | _T_353; // @[LZD.scala 39:25]
  assign _T_355 = {_T_350,_T_354}; // @[Cat.scala 29:58]
  assign _T_356 = _T_348[1]; // @[Shift.scala 12:21]
  assign _T_357 = _T_355[1]; // @[Shift.scala 12:21]
  assign _T_358 = _T_356 | _T_357; // @[LZD.scala 49:16]
  assign _T_359 = ~ _T_357; // @[LZD.scala 49:27]
  assign _T_360 = _T_356 | _T_359; // @[LZD.scala 49:25]
  assign _T_361 = _T_348[0:0]; // @[LZD.scala 49:47]
  assign _T_362 = _T_355[0:0]; // @[LZD.scala 49:59]
  assign _T_363 = _T_356 ? _T_361 : _T_362; // @[LZD.scala 49:35]
  assign _T_365 = {_T_358,_T_360,_T_363}; // @[Cat.scala 29:58]
  assign _T_366 = _T_340[2]; // @[Shift.scala 12:21]
  assign _T_367 = _T_365[2]; // @[Shift.scala 12:21]
  assign _T_368 = _T_366 | _T_367; // @[LZD.scala 49:16]
  assign _T_369 = ~ _T_367; // @[LZD.scala 49:27]
  assign _T_370 = _T_366 | _T_369; // @[LZD.scala 49:25]
  assign _T_371 = _T_340[1:0]; // @[LZD.scala 49:47]
  assign _T_372 = _T_365[1:0]; // @[LZD.scala 49:59]
  assign _T_373 = _T_366 ? _T_371 : _T_372; // @[LZD.scala 49:35]
  assign _T_375 = {_T_368,_T_370,_T_373}; // @[Cat.scala 29:58]
  assign _T_376 = _T_314[7:0]; // @[LZD.scala 44:32]
  assign _T_377 = _T_376[7:4]; // @[LZD.scala 43:32]
  assign _T_378 = _T_377[3:2]; // @[LZD.scala 43:32]
  assign _T_379 = _T_378 != 2'h0; // @[LZD.scala 39:14]
  assign _T_380 = _T_378[1]; // @[LZD.scala 39:21]
  assign _T_381 = _T_378[0]; // @[LZD.scala 39:30]
  assign _T_382 = ~ _T_381; // @[LZD.scala 39:27]
  assign _T_383 = _T_380 | _T_382; // @[LZD.scala 39:25]
  assign _T_384 = {_T_379,_T_383}; // @[Cat.scala 29:58]
  assign _T_385 = _T_377[1:0]; // @[LZD.scala 44:32]
  assign _T_386 = _T_385 != 2'h0; // @[LZD.scala 39:14]
  assign _T_387 = _T_385[1]; // @[LZD.scala 39:21]
  assign _T_388 = _T_385[0]; // @[LZD.scala 39:30]
  assign _T_389 = ~ _T_388; // @[LZD.scala 39:27]
  assign _T_390 = _T_387 | _T_389; // @[LZD.scala 39:25]
  assign _T_391 = {_T_386,_T_390}; // @[Cat.scala 29:58]
  assign _T_392 = _T_384[1]; // @[Shift.scala 12:21]
  assign _T_393 = _T_391[1]; // @[Shift.scala 12:21]
  assign _T_394 = _T_392 | _T_393; // @[LZD.scala 49:16]
  assign _T_395 = ~ _T_393; // @[LZD.scala 49:27]
  assign _T_396 = _T_392 | _T_395; // @[LZD.scala 49:25]
  assign _T_397 = _T_384[0:0]; // @[LZD.scala 49:47]
  assign _T_398 = _T_391[0:0]; // @[LZD.scala 49:59]
  assign _T_399 = _T_392 ? _T_397 : _T_398; // @[LZD.scala 49:35]
  assign _T_401 = {_T_394,_T_396,_T_399}; // @[Cat.scala 29:58]
  assign _T_402 = _T_376[3:0]; // @[LZD.scala 44:32]
  assign _T_403 = _T_402[3:2]; // @[LZD.scala 43:32]
  assign _T_404 = _T_403 != 2'h0; // @[LZD.scala 39:14]
  assign _T_405 = _T_403[1]; // @[LZD.scala 39:21]
  assign _T_406 = _T_403[0]; // @[LZD.scala 39:30]
  assign _T_407 = ~ _T_406; // @[LZD.scala 39:27]
  assign _T_408 = _T_405 | _T_407; // @[LZD.scala 39:25]
  assign _T_409 = {_T_404,_T_408}; // @[Cat.scala 29:58]
  assign _T_410 = _T_402[1:0]; // @[LZD.scala 44:32]
  assign _T_411 = _T_410 != 2'h0; // @[LZD.scala 39:14]
  assign _T_412 = _T_410[1]; // @[LZD.scala 39:21]
  assign _T_413 = _T_410[0]; // @[LZD.scala 39:30]
  assign _T_414 = ~ _T_413; // @[LZD.scala 39:27]
  assign _T_415 = _T_412 | _T_414; // @[LZD.scala 39:25]
  assign _T_416 = {_T_411,_T_415}; // @[Cat.scala 29:58]
  assign _T_417 = _T_409[1]; // @[Shift.scala 12:21]
  assign _T_418 = _T_416[1]; // @[Shift.scala 12:21]
  assign _T_419 = _T_417 | _T_418; // @[LZD.scala 49:16]
  assign _T_420 = ~ _T_418; // @[LZD.scala 49:27]
  assign _T_421 = _T_417 | _T_420; // @[LZD.scala 49:25]
  assign _T_422 = _T_409[0:0]; // @[LZD.scala 49:47]
  assign _T_423 = _T_416[0:0]; // @[LZD.scala 49:59]
  assign _T_424 = _T_417 ? _T_422 : _T_423; // @[LZD.scala 49:35]
  assign _T_426 = {_T_419,_T_421,_T_424}; // @[Cat.scala 29:58]
  assign _T_427 = _T_401[2]; // @[Shift.scala 12:21]
  assign _T_428 = _T_426[2]; // @[Shift.scala 12:21]
  assign _T_429 = _T_427 | _T_428; // @[LZD.scala 49:16]
  assign _T_430 = ~ _T_428; // @[LZD.scala 49:27]
  assign _T_431 = _T_427 | _T_430; // @[LZD.scala 49:25]
  assign _T_432 = _T_401[1:0]; // @[LZD.scala 49:47]
  assign _T_433 = _T_426[1:0]; // @[LZD.scala 49:59]
  assign _T_434 = _T_427 ? _T_432 : _T_433; // @[LZD.scala 49:35]
  assign _T_436 = {_T_429,_T_431,_T_434}; // @[Cat.scala 29:58]
  assign _T_437 = _T_375[3]; // @[Shift.scala 12:21]
  assign _T_438 = _T_436[3]; // @[Shift.scala 12:21]
  assign _T_439 = _T_437 | _T_438; // @[LZD.scala 49:16]
  assign _T_440 = ~ _T_438; // @[LZD.scala 49:27]
  assign _T_441 = _T_437 | _T_440; // @[LZD.scala 49:25]
  assign _T_442 = _T_375[2:0]; // @[LZD.scala 49:47]
  assign _T_443 = _T_436[2:0]; // @[LZD.scala 49:59]
  assign _T_444 = _T_437 ? _T_442 : _T_443; // @[LZD.scala 49:35]
  assign _T_446 = {_T_439,_T_441,_T_444}; // @[Cat.scala 29:58]
  assign _T_447 = _T_313[13:0]; // @[LZD.scala 44:32]
  assign _T_448 = _T_447[13:6]; // @[LZD.scala 43:32]
  assign _T_449 = _T_448[7:4]; // @[LZD.scala 43:32]
  assign _T_450 = _T_449[3:2]; // @[LZD.scala 43:32]
  assign _T_451 = _T_450 != 2'h0; // @[LZD.scala 39:14]
  assign _T_452 = _T_450[1]; // @[LZD.scala 39:21]
  assign _T_453 = _T_450[0]; // @[LZD.scala 39:30]
  assign _T_454 = ~ _T_453; // @[LZD.scala 39:27]
  assign _T_455 = _T_452 | _T_454; // @[LZD.scala 39:25]
  assign _T_456 = {_T_451,_T_455}; // @[Cat.scala 29:58]
  assign _T_457 = _T_449[1:0]; // @[LZD.scala 44:32]
  assign _T_458 = _T_457 != 2'h0; // @[LZD.scala 39:14]
  assign _T_459 = _T_457[1]; // @[LZD.scala 39:21]
  assign _T_460 = _T_457[0]; // @[LZD.scala 39:30]
  assign _T_461 = ~ _T_460; // @[LZD.scala 39:27]
  assign _T_462 = _T_459 | _T_461; // @[LZD.scala 39:25]
  assign _T_463 = {_T_458,_T_462}; // @[Cat.scala 29:58]
  assign _T_464 = _T_456[1]; // @[Shift.scala 12:21]
  assign _T_465 = _T_463[1]; // @[Shift.scala 12:21]
  assign _T_466 = _T_464 | _T_465; // @[LZD.scala 49:16]
  assign _T_467 = ~ _T_465; // @[LZD.scala 49:27]
  assign _T_468 = _T_464 | _T_467; // @[LZD.scala 49:25]
  assign _T_469 = _T_456[0:0]; // @[LZD.scala 49:47]
  assign _T_470 = _T_463[0:0]; // @[LZD.scala 49:59]
  assign _T_471 = _T_464 ? _T_469 : _T_470; // @[LZD.scala 49:35]
  assign _T_473 = {_T_466,_T_468,_T_471}; // @[Cat.scala 29:58]
  assign _T_474 = _T_448[3:0]; // @[LZD.scala 44:32]
  assign _T_475 = _T_474[3:2]; // @[LZD.scala 43:32]
  assign _T_476 = _T_475 != 2'h0; // @[LZD.scala 39:14]
  assign _T_477 = _T_475[1]; // @[LZD.scala 39:21]
  assign _T_478 = _T_475[0]; // @[LZD.scala 39:30]
  assign _T_479 = ~ _T_478; // @[LZD.scala 39:27]
  assign _T_480 = _T_477 | _T_479; // @[LZD.scala 39:25]
  assign _T_481 = {_T_476,_T_480}; // @[Cat.scala 29:58]
  assign _T_482 = _T_474[1:0]; // @[LZD.scala 44:32]
  assign _T_483 = _T_482 != 2'h0; // @[LZD.scala 39:14]
  assign _T_484 = _T_482[1]; // @[LZD.scala 39:21]
  assign _T_485 = _T_482[0]; // @[LZD.scala 39:30]
  assign _T_486 = ~ _T_485; // @[LZD.scala 39:27]
  assign _T_487 = _T_484 | _T_486; // @[LZD.scala 39:25]
  assign _T_488 = {_T_483,_T_487}; // @[Cat.scala 29:58]
  assign _T_489 = _T_481[1]; // @[Shift.scala 12:21]
  assign _T_490 = _T_488[1]; // @[Shift.scala 12:21]
  assign _T_491 = _T_489 | _T_490; // @[LZD.scala 49:16]
  assign _T_492 = ~ _T_490; // @[LZD.scala 49:27]
  assign _T_493 = _T_489 | _T_492; // @[LZD.scala 49:25]
  assign _T_494 = _T_481[0:0]; // @[LZD.scala 49:47]
  assign _T_495 = _T_488[0:0]; // @[LZD.scala 49:59]
  assign _T_496 = _T_489 ? _T_494 : _T_495; // @[LZD.scala 49:35]
  assign _T_498 = {_T_491,_T_493,_T_496}; // @[Cat.scala 29:58]
  assign _T_499 = _T_473[2]; // @[Shift.scala 12:21]
  assign _T_500 = _T_498[2]; // @[Shift.scala 12:21]
  assign _T_501 = _T_499 | _T_500; // @[LZD.scala 49:16]
  assign _T_502 = ~ _T_500; // @[LZD.scala 49:27]
  assign _T_503 = _T_499 | _T_502; // @[LZD.scala 49:25]
  assign _T_504 = _T_473[1:0]; // @[LZD.scala 49:47]
  assign _T_505 = _T_498[1:0]; // @[LZD.scala 49:59]
  assign _T_506 = _T_499 ? _T_504 : _T_505; // @[LZD.scala 49:35]
  assign _T_508 = {_T_501,_T_503,_T_506}; // @[Cat.scala 29:58]
  assign _T_509 = _T_447[5:0]; // @[LZD.scala 44:32]
  assign _T_510 = _T_509[5:2]; // @[LZD.scala 43:32]
  assign _T_511 = _T_510[3:2]; // @[LZD.scala 43:32]
  assign _T_512 = _T_511 != 2'h0; // @[LZD.scala 39:14]
  assign _T_513 = _T_511[1]; // @[LZD.scala 39:21]
  assign _T_514 = _T_511[0]; // @[LZD.scala 39:30]
  assign _T_515 = ~ _T_514; // @[LZD.scala 39:27]
  assign _T_516 = _T_513 | _T_515; // @[LZD.scala 39:25]
  assign _T_517 = {_T_512,_T_516}; // @[Cat.scala 29:58]
  assign _T_518 = _T_510[1:0]; // @[LZD.scala 44:32]
  assign _T_519 = _T_518 != 2'h0; // @[LZD.scala 39:14]
  assign _T_520 = _T_518[1]; // @[LZD.scala 39:21]
  assign _T_521 = _T_518[0]; // @[LZD.scala 39:30]
  assign _T_522 = ~ _T_521; // @[LZD.scala 39:27]
  assign _T_523 = _T_520 | _T_522; // @[LZD.scala 39:25]
  assign _T_524 = {_T_519,_T_523}; // @[Cat.scala 29:58]
  assign _T_525 = _T_517[1]; // @[Shift.scala 12:21]
  assign _T_526 = _T_524[1]; // @[Shift.scala 12:21]
  assign _T_527 = _T_525 | _T_526; // @[LZD.scala 49:16]
  assign _T_528 = ~ _T_526; // @[LZD.scala 49:27]
  assign _T_529 = _T_525 | _T_528; // @[LZD.scala 49:25]
  assign _T_530 = _T_517[0:0]; // @[LZD.scala 49:47]
  assign _T_531 = _T_524[0:0]; // @[LZD.scala 49:59]
  assign _T_532 = _T_525 ? _T_530 : _T_531; // @[LZD.scala 49:35]
  assign _T_534 = {_T_527,_T_529,_T_532}; // @[Cat.scala 29:58]
  assign _T_535 = _T_509[1:0]; // @[LZD.scala 44:32]
  assign _T_536 = _T_535 != 2'h0; // @[LZD.scala 39:14]
  assign _T_537 = _T_535[1]; // @[LZD.scala 39:21]
  assign _T_538 = _T_535[0]; // @[LZD.scala 39:30]
  assign _T_539 = ~ _T_538; // @[LZD.scala 39:27]
  assign _T_540 = _T_537 | _T_539; // @[LZD.scala 39:25]
  assign _T_541 = {_T_536,_T_540}; // @[Cat.scala 29:58]
  assign _T_542 = _T_534[2]; // @[Shift.scala 12:21]
  assign _T_544 = _T_534[1:0]; // @[LZD.scala 55:32]
  assign _T_545 = _T_542 ? _T_544 : _T_541; // @[LZD.scala 55:20]
  assign _T_546 = {_T_542,_T_545}; // @[Cat.scala 29:58]
  assign _T_547 = _T_508[3]; // @[Shift.scala 12:21]
  assign _T_549 = _T_508[2:0]; // @[LZD.scala 55:32]
  assign _T_550 = _T_547 ? _T_549 : _T_546; // @[LZD.scala 55:20]
  assign _T_551 = {_T_547,_T_550}; // @[Cat.scala 29:58]
  assign _T_552 = _T_446[4]; // @[Shift.scala 12:21]
  assign _T_554 = _T_446[3:0]; // @[LZD.scala 55:32]
  assign _T_555 = _T_552 ? _T_554 : _T_551; // @[LZD.scala 55:20]
  assign _T_556 = {_T_552,_T_555}; // @[Cat.scala 29:58]
  assign _T_557 = ~ _T_556; // @[convert.scala 21:22]
  assign _T_558 = io_B[28:0]; // @[convert.scala 22:36]
  assign _T_559 = _T_557 < 5'h1d; // @[Shift.scala 16:24]
  assign _T_561 = _T_557[4]; // @[Shift.scala 12:21]
  assign _T_562 = _T_558[12:0]; // @[Shift.scala 64:52]
  assign _T_564 = {_T_562,16'h0}; // @[Cat.scala 29:58]
  assign _T_565 = _T_561 ? _T_564 : _T_558; // @[Shift.scala 64:27]
  assign _T_566 = _T_557[3:0]; // @[Shift.scala 66:70]
  assign _T_567 = _T_566[3]; // @[Shift.scala 12:21]
  assign _T_568 = _T_565[20:0]; // @[Shift.scala 64:52]
  assign _T_570 = {_T_568,8'h0}; // @[Cat.scala 29:58]
  assign _T_571 = _T_567 ? _T_570 : _T_565; // @[Shift.scala 64:27]
  assign _T_572 = _T_566[2:0]; // @[Shift.scala 66:70]
  assign _T_573 = _T_572[2]; // @[Shift.scala 12:21]
  assign _T_574 = _T_571[24:0]; // @[Shift.scala 64:52]
  assign _T_576 = {_T_574,4'h0}; // @[Cat.scala 29:58]
  assign _T_577 = _T_573 ? _T_576 : _T_571; // @[Shift.scala 64:27]
  assign _T_578 = _T_572[1:0]; // @[Shift.scala 66:70]
  assign _T_579 = _T_578[1]; // @[Shift.scala 12:21]
  assign _T_580 = _T_577[26:0]; // @[Shift.scala 64:52]
  assign _T_582 = {_T_580,2'h0}; // @[Cat.scala 29:58]
  assign _T_583 = _T_579 ? _T_582 : _T_577; // @[Shift.scala 64:27]
  assign _T_584 = _T_578[0:0]; // @[Shift.scala 66:70]
  assign _T_586 = _T_583[27:0]; // @[Shift.scala 64:52]
  assign _T_587 = {_T_586,1'h0}; // @[Cat.scala 29:58]
  assign _T_588 = _T_584 ? _T_587 : _T_583; // @[Shift.scala 64:27]
  assign _T_589 = _T_559 ? _T_588 : 29'h0; // @[Shift.scala 16:10]
  assign _T_590 = _T_589[28:28]; // @[convert.scala 23:34]
  assign decB_fraction = _T_589[27:0]; // @[convert.scala 24:34]
  assign _T_592 = _T_310 == 1'h0; // @[convert.scala 25:26]
  assign _T_594 = _T_310 ? _T_557 : _T_556; // @[convert.scala 25:42]
  assign _T_597 = ~ _T_590; // @[convert.scala 26:67]
  assign _T_598 = _T_308 ? _T_597 : _T_590; // @[convert.scala 26:51]
  assign _T_599 = {_T_592,_T_594,_T_598}; // @[Cat.scala 29:58]
  assign _T_601 = io_B[30:0]; // @[convert.scala 29:56]
  assign _T_602 = _T_601 != 31'h0; // @[convert.scala 29:60]
  assign _T_603 = ~ _T_602; // @[convert.scala 29:41]
  assign decB_isNaR = _T_308 & _T_603; // @[convert.scala 29:39]
  assign _T_606 = _T_308 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_606 & _T_603; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_599); // @[convert.scala 32:24]
  assign _T_615 = _T_1 ? 3'h7 : 3'h0; // @[Bitwise.scala 71:12]
  assign _T_616 = ~ _T_1; // @[PositDivisionSqrt.scala 80:40]
  assign sigA_S = {_T_615,_T_616,decA_fraction,3'h0}; // @[Cat.scala 29:58]
  assign _T_619 = ~ _T_308; // @[PositDivisionSqrt.scala 82:31]
  assign sigB_S = {_T_308,_T_619,decB_fraction,5'h0}; // @[Cat.scala 29:58]
  assign _T_622 = decA_isNaR == 1'h0; // @[PositDivisionSqrt.scala 85:25]
  assign invalidSqrt = _T_622 & _T_1; // @[PositDivisionSqrt.scala 85:37]
  assign _T_623 = decA_isNaR | invalidSqrt; // @[PositDivisionSqrt.scala 88:42]
  assign _T_624 = decA_isNaR | decB_isNaR; // @[PositDivisionSqrt.scala 89:42]
  assign _T_625 = _T_624 | decB_isZero; // @[PositDivisionSqrt.scala 89:56]
  assign _T_626 = decB_isZero == 1'h0; // @[PositDivisionSqrt.scala 94:46]
  assign _T_627 = decA_isZero & _T_626; // @[PositDivisionSqrt.scala 94:43]
  assign _T_628 = decB_isNaR == 1'h0; // @[PositDivisionSqrt.scala 94:62]
  assign _T_629 = _T_627 & _T_628; // @[PositDivisionSqrt.scala 94:59]
  assign specialCaseA_S = decA_isNaR | decA_isZero; // @[PositDivisionSqrt.scala 97:38]
  assign specialCaseB_S = decB_isNaR | decB_isZero; // @[PositDivisionSqrt.scala 98:38]
  assign _T_630 = specialCaseA_S == 1'h0; // @[PositDivisionSqrt.scala 99:27]
  assign _T_631 = specialCaseB_S == 1'h0; // @[PositDivisionSqrt.scala 99:46]
  assign normalCase_S_div = _T_630 & _T_631; // @[PositDivisionSqrt.scala 99:43]
  assign normalCase_S_sqrt = _T_630 & _T_299; // @[PositDivisionSqrt.scala 100:43]
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div; // @[PositDivisionSqrt.scala 101:30]
  assign sExpQuot_S_div = $signed(decA_scale) - $signed(decB_scale); // @[PositDivisionSqrt.scala 103:38]
  assign _T_634 = decA_scale[0]; // @[PositDivisionSqrt.scala 104:50]
  assign oddSqrt_S = io_sqrtOp & _T_634; // @[PositDivisionSqrt.scala 104:37]
  assign idle = cycleNum == 6'h0; // @[PositDivisionSqrt.scala 109:39]
  assign ready = cycleNum <= 6'h1; // @[PositDivisionSqrt.scala 110:39]
  assign entering = ready & io_inValid; // @[PositDivisionSqrt.scala 111:35]
  assign entering_normalCase = entering & normalCase_S; // @[PositDivisionSqrt.scala 112:38]
  assign _T_635 = sigX_Z[34]; // @[PositDivisionSqrt.scala 113:35]
  assign _T_636 = sigX_Z[32]; // @[PositDivisionSqrt.scala 113:58]
  assign scaleNotChange = _T_635 ^ _T_636; // @[PositDivisionSqrt.scala 113:50]
  assign _T_637 = cycleNum == 6'h3; // @[PositDivisionSqrt.scala 114:39]
  assign skipCycle2 = _T_637 & scaleNotChange; // @[PositDivisionSqrt.scala 114:48]
  assign _T_638 = idle == 1'h0; // @[PositDivisionSqrt.scala 116:8]
  assign _T_639 = _T_638 | io_inValid; // @[PositDivisionSqrt.scala 116:14]
  assign _T_640 = normalCase_S == 1'h0; // @[PositDivisionSqrt.scala 117:32]
  assign _T_641 = entering & _T_640; // @[PositDivisionSqrt.scala 117:30]
  assign _T_643 = io_sqrtOp ? 6'h21 : 6'h23; // @[PositDivisionSqrt.scala 119:26]
  assign _T_644 = entering_normalCase ? _T_643 : 6'h0; // @[PositDivisionSqrt.scala 118:20]
  assign _GEN_9 = {{5'd0}, _T_641}; // @[PositDivisionSqrt.scala 117:64]
  assign _T_645 = _GEN_9 | _T_644; // @[PositDivisionSqrt.scala 117:64]
  assign _T_647 = skipCycle2 == 1'h0; // @[PositDivisionSqrt.scala 123:30]
  assign _T_648 = _T_638 & _T_647; // @[PositDivisionSqrt.scala 123:27]
  assign _T_650 = cycleNum - 6'h1; // @[PositDivisionSqrt.scala 123:52]
  assign _T_651 = _T_648 ? _T_650 : 6'h0; // @[PositDivisionSqrt.scala 123:20]
  assign _T_652 = _T_645 | _T_651; // @[PositDivisionSqrt.scala 122:64]
  assign _T_654 = _T_638 & skipCycle2; // @[PositDivisionSqrt.scala 124:27]
  assign _GEN_10 = {{5'd0}, _T_654}; // @[PositDivisionSqrt.scala 123:64]
  assign _T_656 = _T_652 | _GEN_10; // @[PositDivisionSqrt.scala 123:64]
  assign _T_657 = decA_scale[6:1]; // @[PositDivisionSqrt.scala 134:42]
  assign _T_659 = io_sqrtOp == 1'h0; // @[PositDivisionSqrt.scala 137:31]
  assign _T_660 = entering_normalCase & _T_659; // @[PositDivisionSqrt.scala 137:28]
  assign _T_661 = 64'h1 << cycleNum; // @[PositDivisionSqrt.scala 146:22]
  assign _T_662 = _T_661[63:2]; // @[PositDivisionSqrt.scala 146:35]
  assign _T_663 = oddSqrt_S == 1'h0; // @[PositDivisionSqrt.scala 148:26]
  assign _T_664 = ready & _T_663; // @[PositDivisionSqrt.scala 148:23]
  assign _T_665 = _T_664 ? sigA_S : 35'h0; // @[PositDivisionSqrt.scala 148:16]
  assign _T_666 = ready & oddSqrt_S; // @[PositDivisionSqrt.scala 149:23]
  assign _T_667 = {sigA_S, 1'h0}; // @[PositDivisionSqrt.scala 149:46]
  assign _T_668 = _T_667[34:0]; // @[PositDivisionSqrt.scala 149:56]
  assign _T_669 = _T_666 ? _T_668 : 35'h0; // @[PositDivisionSqrt.scala 149:16]
  assign _T_670 = _T_665 | _T_669; // @[PositDivisionSqrt.scala 148:66]
  assign _T_671 = ready == 1'h0; // @[PositDivisionSqrt.scala 150:17]
  assign _T_672 = _T_671 ? rem_Z : 35'h0; // @[PositDivisionSqrt.scala 150:16]
  assign rem = _T_670 | _T_672; // @[PositDivisionSqrt.scala 149:66]
  assign _T_674 = ready & _T_659; // @[PositDivisionSqrt.scala 152:29]
  assign _T_675 = _T_674 ? sigB_S : 35'h0; // @[PositDivisionSqrt.scala 152:22]
  assign _T_676 = ready & io_sqrtOp; // @[PositDivisionSqrt.scala 153:29]
  assign _T_677 = _T_676 ? 32'h80000000 : 32'h0; // @[PositDivisionSqrt.scala 153:22]
  assign _GEN_11 = {{3'd0}, _T_677}; // @[PositDivisionSqrt.scala 152:93]
  assign _T_678 = _T_675 | _GEN_11; // @[PositDivisionSqrt.scala 152:93]
  assign _T_680 = sqrtOp_Z == 1'h0; // @[PositDivisionSqrt.scala 154:33]
  assign _T_681 = _T_671 & _T_680; // @[PositDivisionSqrt.scala 154:30]
  assign _T_682 = ~ signB_Z; // @[PositDivisionSqrt.scala 154:57]
  assign _T_685 = {signB_Z,_T_682,fractB_Z,5'h0}; // @[Cat.scala 29:58]
  assign _T_686 = _T_681 ? _T_685 : 35'h0; // @[PositDivisionSqrt.scala 154:22]
  assign _T_687 = _T_678 | _T_686; // @[PositDivisionSqrt.scala 153:93]
  assign _T_689 = _T_671 & sqrtOp_Z; // @[PositDivisionSqrt.scala 155:30]
  assign _T_690 = rem[34:34]; // @[PositDivisionSqrt.scala 156:83]
  assign _T_692 = _T_690 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 71:12]
  assign bitMask = _T_662[33:0]; // @[PositDivisionSqrt.scala 145:21 PositDivisionSqrt.scala 146:14]
  assign _GEN_12 = {{3'd0}, _T_692}; // @[PositDivisionSqrt.scala 156:53]
  assign _T_693 = bitMask & _GEN_12; // @[PositDivisionSqrt.scala 156:53]
  assign _GEN_13 = {{1'd0}, _T_693}; // @[PositDivisionSqrt.scala 155:51]
  assign _T_694 = sigX_Z | _GEN_13; // @[PositDivisionSqrt.scala 155:51]
  assign _T_695 = bitMask[33:1]; // @[PositDivisionSqrt.scala 157:53]
  assign _GEN_14 = {{2'd0}, _T_695}; // @[PositDivisionSqrt.scala 156:89]
  assign _T_696 = _T_694 | _GEN_14; // @[PositDivisionSqrt.scala 156:89]
  assign _T_697 = _T_689 ? _T_696 : 35'h0; // @[PositDivisionSqrt.scala 155:22]
  assign trialTerm = _T_687 | _T_697; // @[PositDivisionSqrt.scala 154:93]
  assign _T_699 = trialTerm[34:34]; // @[PositDivisionSqrt.scala 162:56]
  assign _T_700 = _T_690 ^ _T_699; // @[PositDivisionSqrt.scala 162:40]
  assign _T_703 = rem + trialTerm; // @[PositDivisionSqrt.scala 163:97]
  assign _T_705 = rem - trialTerm; // @[PositDivisionSqrt.scala 164:97]
  assign _T_706 = _T_700 ? _T_703 : _T_705; // @[PositDivisionSqrt.scala 161:92]
  assign _T_711 = {rem, 1'h0}; // @[PositDivisionSqrt.scala 168:98]
  assign _T_712 = _T_711[34:0]; // @[PositDivisionSqrt.scala 168:108]
  assign _T_714 = _T_712 + trialTerm; // @[PositDivisionSqrt.scala 168:112]
  assign _T_718 = _T_712 - trialTerm; // @[PositDivisionSqrt.scala 169:112]
  assign _T_719 = _T_700 ? _T_714 : _T_718; // @[PositDivisionSqrt.scala 166:26]
  assign trialRem = ready ? _T_706 : _T_719; // @[PositDivisionSqrt.scala 159:27]
  assign _T_720 = trialRem != 35'h0; // @[PositDivisionSqrt.scala 173:35]
  assign trIsZero = _T_720 == 1'h0; // @[PositDivisionSqrt.scala 173:25]
  assign _T_721 = rem != 35'h0; // @[PositDivisionSqrt.scala 174:30]
  assign remIsZero = _T_721 == 1'h0; // @[PositDivisionSqrt.scala 174:25]
  assign _T_723 = trialRem[34:34]; // @[PositDivisionSqrt.scala 176:64]
  assign _T_724 = _T_699 ^ _T_723; // @[PositDivisionSqrt.scala 176:49]
  assign _T_725 = ~ _T_724; // @[PositDivisionSqrt.scala 176:29]
  assign _T_726 = sigX_Z[34:34]; // @[PositDivisionSqrt.scala 178:61]
  assign _T_727 = ~ _T_726; // @[PositDivisionSqrt.scala 178:49]
  assign _T_729 = remIsZero ? _T_726 : _T_725; // @[Mux.scala 87:16]
  assign newBit = trIsZero ? _T_727 : _T_729; // @[Mux.scala 87:16]
  assign _T_730 = cycleNum > 6'h2; // @[PositDivisionSqrt.scala 183:41]
  assign _T_731 = remIsZero == 1'h0; // @[PositDivisionSqrt.scala 183:51]
  assign _T_732 = _T_730 & _T_731; // @[PositDivisionSqrt.scala 183:48]
  assign _T_733 = entering_normalCase | _T_732; // @[PositDivisionSqrt.scala 183:28]
  assign _T_736 = _T_671 & newBit; // @[PositDivisionSqrt.scala 187:39]
  assign _T_737 = entering_normalCase | _T_736; // @[PositDivisionSqrt.scala 187:28]
  assign _T_740 = {newBit, 34'h0}; // @[PositDivisionSqrt.scala 188:47]
  assign _T_741 = _T_674 ? _T_740 : 35'h0; // @[PositDivisionSqrt.scala 188:18]
  assign _T_743 = _T_676 ? 33'h100000000 : 33'h0; // @[PositDivisionSqrt.scala 189:18]
  assign _GEN_15 = {{2'd0}, _T_743}; // @[PositDivisionSqrt.scala 188:78]
  assign _T_744 = _T_741 | _GEN_15; // @[PositDivisionSqrt.scala 188:78]
  assign _GEN_16 = {{1'd0}, bitMask}; // @[PositDivisionSqrt.scala 190:47]
  assign _T_746 = sigX_Z | _GEN_16; // @[PositDivisionSqrt.scala 190:47]
  assign _T_747 = _T_671 ? _T_746 : 35'h0; // @[PositDivisionSqrt.scala 190:18]
  assign _T_748 = _T_744 | _T_747; // @[PositDivisionSqrt.scala 189:78]
  assign _T_750 = {_T_726, 1'h0}; // @[PositDivisionSqrt.scala 196:53]
  assign sigXBias = scaleNotChange ? _T_750 : {{1'd0}, _T_726}; // @[PositDivisionSqrt.scala 196:21]
  assign _GEN_17 = {{33'd0}, sigXBias}; // @[PositDivisionSqrt.scala 197:25]
  assign realSigX = sigX_Z + _GEN_17; // @[PositDivisionSqrt.scala 197:25]
  assign _T_753 = realSigX[31:4]; // @[PositDivisionSqrt.scala 200:97]
  assign _T_754 = realSigX[30:3]; // @[PositDivisionSqrt.scala 201:97]
  assign realFrac = scaleNotChange ? _T_753 : _T_754; // @[PositDivisionSqrt.scala 198:21]
  assign _T_755 = realSigX[34]; // @[PositDivisionSqrt.scala 205:33]
  assign _T_756 = realSigX[32]; // @[PositDivisionSqrt.scala 205:58]
  assign _T_757 = _T_755 ^ _T_756; // @[PositDivisionSqrt.scala 205:48]
  assign scaleNeedSub = ~ _T_757; // @[PositDivisionSqrt.scala 205:23]
  assign _T_759 = realSigX[31]; // @[PositDivisionSqrt.scala 206:56]
  assign notNeedSubTwo = _T_755 ^ _T_759; // @[PositDivisionSqrt.scala 206:46]
  assign scaleSubOne = scaleNeedSub & notNeedSubTwo; // @[PositDivisionSqrt.scala 207:36]
  assign _T_760 = ~ notNeedSubTwo; // @[PositDivisionSqrt.scala 208:38]
  assign scaleSubTwo = scaleNeedSub & _T_760; // @[PositDivisionSqrt.scala 208:36]
  assign _T_761 = {scaleSubTwo,scaleSubOne}; // @[Cat.scala 29:58]
  assign _T_762 = {1'b0,$signed(_T_761)}; // @[PositDivisionSqrt.scala 209:63]
  assign _GEN_18 = {{5{_T_762[2]}},_T_762}; // @[PositDivisionSqrt.scala 209:31]
  assign _T_764 = $signed(scale_Z) - $signed(_GEN_18); // @[PositDivisionSqrt.scala 209:31]
  assign realExp = $signed(_T_764); // @[PositDivisionSqrt.scala 209:31]
  assign underflow = $signed(realExp) < $signed(-8'sh3d); // @[PositDivisionSqrt.scala 210:31]
  assign overflow = $signed(realExp) > $signed(8'sh3c); // @[PositDivisionSqrt.scala 211:31]
  assign decQ_sign = realSigX[34:34]; // @[PositDivisionSqrt.scala 215:33]
  assign _T_766 = underflow ? $signed(-8'sh3d) : $signed(realExp); // @[Mux.scala 87:16]
  assign _T_767 = overflow ? $signed(8'sh3c) : $signed(_T_766); // @[Mux.scala 87:16]
  assign _T_768 = realSigX[3:1]; // @[PositDivisionSqrt.scala 224:48]
  assign _T_769 = realSigX[2:0]; // @[PositDivisionSqrt.scala 224:64]
  assign decQ_grs = scaleNotChange ? _T_768 : _T_769; // @[PositDivisionSqrt.scala 224:23]
  assign outValid = cycleNum == 6'h1; // @[PositDivisionSqrt.scala 229:28]
  assign _GEN_19 = _T_767[6:0]; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign decQ_scale = $signed(_GEN_19); // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign _T_775 = decQ_scale[0]; // @[convert.scala 46:61]
  assign _T_776 = ~ _T_775; // @[convert.scala 46:52]
  assign _T_778 = decQ_sign ? _T_776 : _T_775; // @[convert.scala 46:42]
  assign _T_779 = decQ_scale[6:1]; // @[convert.scala 48:34]
  assign _T_780 = _T_779[5:5]; // @[convert.scala 49:36]
  assign _T_782 = ~ _T_779; // @[convert.scala 50:36]
  assign _T_783 = $signed(_T_782); // @[convert.scala 50:36]
  assign _T_784 = _T_780 ? $signed(_T_783) : $signed(_T_779); // @[convert.scala 50:28]
  assign _T_785 = _T_780 ^ decQ_sign; // @[convert.scala 51:31]
  assign _T_786 = ~ _T_785; // @[convert.scala 52:43]
  assign _T_790 = {_T_786,_T_785,_T_778,realFrac,decQ_grs}; // @[Cat.scala 29:58]
  assign _T_791 = $unsigned(_T_784); // @[Shift.scala 39:17]
  assign _T_792 = _T_791 < 6'h22; // @[Shift.scala 39:24]
  assign _T_794 = _T_790[33:32]; // @[Shift.scala 90:30]
  assign _T_795 = _T_790[31:0]; // @[Shift.scala 90:48]
  assign _T_796 = _T_795 != 32'h0; // @[Shift.scala 90:57]
  assign _GEN_20 = {{1'd0}, _T_796}; // @[Shift.scala 90:39]
  assign _T_797 = _T_794 | _GEN_20; // @[Shift.scala 90:39]
  assign _T_798 = _T_791[5]; // @[Shift.scala 12:21]
  assign _T_799 = _T_790[33]; // @[Shift.scala 12:21]
  assign _T_801 = _T_799 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 71:12]
  assign _T_802 = {_T_801,_T_797}; // @[Cat.scala 29:58]
  assign _T_803 = _T_798 ? _T_802 : _T_790; // @[Shift.scala 91:22]
  assign _T_804 = _T_791[4:0]; // @[Shift.scala 92:77]
  assign _T_805 = _T_803[33:16]; // @[Shift.scala 90:30]
  assign _T_806 = _T_803[15:0]; // @[Shift.scala 90:48]
  assign _T_807 = _T_806 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_21 = {{17'd0}, _T_807}; // @[Shift.scala 90:39]
  assign _T_808 = _T_805 | _GEN_21; // @[Shift.scala 90:39]
  assign _T_809 = _T_804[4]; // @[Shift.scala 12:21]
  assign _T_810 = _T_803[33]; // @[Shift.scala 12:21]
  assign _T_812 = _T_810 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_813 = {_T_812,_T_808}; // @[Cat.scala 29:58]
  assign _T_814 = _T_809 ? _T_813 : _T_803; // @[Shift.scala 91:22]
  assign _T_815 = _T_804[3:0]; // @[Shift.scala 92:77]
  assign _T_816 = _T_814[33:8]; // @[Shift.scala 90:30]
  assign _T_817 = _T_814[7:0]; // @[Shift.scala 90:48]
  assign _T_818 = _T_817 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_22 = {{25'd0}, _T_818}; // @[Shift.scala 90:39]
  assign _T_819 = _T_816 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_820 = _T_815[3]; // @[Shift.scala 12:21]
  assign _T_821 = _T_814[33]; // @[Shift.scala 12:21]
  assign _T_823 = _T_821 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_824 = {_T_823,_T_819}; // @[Cat.scala 29:58]
  assign _T_825 = _T_820 ? _T_824 : _T_814; // @[Shift.scala 91:22]
  assign _T_826 = _T_815[2:0]; // @[Shift.scala 92:77]
  assign _T_827 = _T_825[33:4]; // @[Shift.scala 90:30]
  assign _T_828 = _T_825[3:0]; // @[Shift.scala 90:48]
  assign _T_829 = _T_828 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_23 = {{29'd0}, _T_829}; // @[Shift.scala 90:39]
  assign _T_830 = _T_827 | _GEN_23; // @[Shift.scala 90:39]
  assign _T_831 = _T_826[2]; // @[Shift.scala 12:21]
  assign _T_832 = _T_825[33]; // @[Shift.scala 12:21]
  assign _T_834 = _T_832 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_835 = {_T_834,_T_830}; // @[Cat.scala 29:58]
  assign _T_836 = _T_831 ? _T_835 : _T_825; // @[Shift.scala 91:22]
  assign _T_837 = _T_826[1:0]; // @[Shift.scala 92:77]
  assign _T_838 = _T_836[33:2]; // @[Shift.scala 90:30]
  assign _T_839 = _T_836[1:0]; // @[Shift.scala 90:48]
  assign _T_840 = _T_839 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_24 = {{31'd0}, _T_840}; // @[Shift.scala 90:39]
  assign _T_841 = _T_838 | _GEN_24; // @[Shift.scala 90:39]
  assign _T_842 = _T_837[1]; // @[Shift.scala 12:21]
  assign _T_843 = _T_836[33]; // @[Shift.scala 12:21]
  assign _T_845 = _T_843 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_846 = {_T_845,_T_841}; // @[Cat.scala 29:58]
  assign _T_847 = _T_842 ? _T_846 : _T_836; // @[Shift.scala 91:22]
  assign _T_848 = _T_837[0:0]; // @[Shift.scala 92:77]
  assign _T_849 = _T_847[33:1]; // @[Shift.scala 90:30]
  assign _T_850 = _T_847[0:0]; // @[Shift.scala 90:48]
  assign _GEN_25 = {{32'd0}, _T_850}; // @[Shift.scala 90:39]
  assign _T_852 = _T_849 | _GEN_25; // @[Shift.scala 90:39]
  assign _T_854 = _T_847[33]; // @[Shift.scala 12:21]
  assign _T_855 = {_T_854,_T_852}; // @[Cat.scala 29:58]
  assign _T_856 = _T_848 ? _T_855 : _T_847; // @[Shift.scala 91:22]
  assign _T_859 = _T_799 ? 34'h3ffffffff : 34'h0; // @[Bitwise.scala 71:12]
  assign _T_860 = _T_792 ? _T_856 : _T_859; // @[Shift.scala 39:10]
  assign _T_861 = _T_860[3]; // @[convert.scala 55:31]
  assign _T_862 = _T_860[2]; // @[convert.scala 56:31]
  assign _T_863 = _T_860[1]; // @[convert.scala 57:31]
  assign _T_864 = _T_860[0]; // @[convert.scala 58:31]
  assign _T_865 = _T_860[33:3]; // @[convert.scala 59:69]
  assign _T_866 = _T_865 != 31'h0; // @[convert.scala 59:81]
  assign _T_867 = ~ _T_866; // @[convert.scala 59:50]
  assign _T_869 = _T_865 == 31'h7fffffff; // @[convert.scala 60:81]
  assign _T_870 = _T_861 | _T_863; // @[convert.scala 61:44]
  assign _T_871 = _T_870 | _T_864; // @[convert.scala 61:52]
  assign _T_872 = _T_862 & _T_871; // @[convert.scala 61:36]
  assign _T_873 = ~ _T_869; // @[convert.scala 62:63]
  assign _T_874 = _T_873 & _T_872; // @[convert.scala 62:103]
  assign _T_875 = _T_867 | _T_874; // @[convert.scala 62:60]
  assign _GEN_26 = {{30'd0}, _T_875}; // @[convert.scala 63:56]
  assign _T_878 = _T_865 + _GEN_26; // @[convert.scala 63:56]
  assign _T_879 = {decQ_sign,_T_878}; // @[Cat.scala 29:58]
  assign _T_881 = isZero_Z ? 32'h0 : _T_879; // @[Mux.scala 87:16]
  assign io_inReady = cycleNum <= 6'h1; // @[PositDivisionSqrt.scala 231:17]
  assign io_diviValid = outValid & _T_680; // @[PositDivisionSqrt.scala 232:17]
  assign io_sqrtValid = outValid & sqrtOp_Z; // @[PositDivisionSqrt.scala 233:17]
  assign io_invalidExc = isNaR_Z; // @[PositDivisionSqrt.scala 234:17]
  assign io_Q = isNaR_Z ? 32'h80000000 : _T_881; // @[PositDivisionSqrt.scala 235:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleNum = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sqrtOp_Z = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  isNaR_Z = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  isZero_Z = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  scale_Z = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  signB_Z = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fractB_Z = _RAND_6[27:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{`RANDOM}};
  rem_Z = _RAND_7[34:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{`RANDOM}};
  sigX_Z = _RAND_8[34:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      cycleNum <= 6'h0;
    end else begin
      if (_T_639) begin
        cycleNum <= _T_656;
      end
    end
    if (entering) begin
      sqrtOp_Z <= io_sqrtOp;
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isNaR_Z <= _T_623;
      end else begin
        isNaR_Z <= _T_625;
      end
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isZero_Z <= decA_isZero;
      end else begin
        isZero_Z <= _T_629;
      end
    end
    if (entering_normalCase) begin
      if (io_sqrtOp) begin
        scale_Z <= {{2{_T_657[5]}},_T_657};
      end else begin
        scale_Z <= sExpQuot_S_div;
      end
    end
    if (_T_660) begin
      signB_Z <= _T_308;
    end
    if (_T_660) begin
      fractB_Z <= decB_fraction;
    end
    if (_T_733) begin
      if (ready) begin
        if (_T_700) begin
          rem_Z <= _T_703;
        end else begin
          rem_Z <= _T_705;
        end
      end else begin
        if (_T_700) begin
          rem_Z <= _T_714;
        end else begin
          rem_Z <= _T_718;
        end
      end
    end
    if (_T_737) begin
      sigX_Z <= _T_748;
    end
  end
endmodule
