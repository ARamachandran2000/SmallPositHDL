module PositAdder16_3(
  input         clock,
  input         reset,
  input  [15:0] io_A,
  input  [15:0] io_B,
  output [15:0] io_S
);
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [13:0] _T_4; // @[convert.scala 19:24]
  wire [13:0] _T_5; // @[convert.scala 19:43]
  wire [13:0] _T_6; // @[convert.scala 19:39]
  wire [7:0] _T_7; // @[LZD.scala 43:32]
  wire [3:0] _T_8; // @[LZD.scala 43:32]
  wire [1:0] _T_9; // @[LZD.scala 43:32]
  wire  _T_10; // @[LZD.scala 39:14]
  wire  _T_11; // @[LZD.scala 39:21]
  wire  _T_12; // @[LZD.scala 39:30]
  wire  _T_13; // @[LZD.scala 39:27]
  wire  _T_14; // @[LZD.scala 39:25]
  wire [1:0] _T_15; // @[Cat.scala 29:58]
  wire [1:0] _T_16; // @[LZD.scala 44:32]
  wire  _T_17; // @[LZD.scala 39:14]
  wire  _T_18; // @[LZD.scala 39:21]
  wire  _T_19; // @[LZD.scala 39:30]
  wire  _T_20; // @[LZD.scala 39:27]
  wire  _T_21; // @[LZD.scala 39:25]
  wire [1:0] _T_22; // @[Cat.scala 29:58]
  wire  _T_23; // @[Shift.scala 12:21]
  wire  _T_24; // @[Shift.scala 12:21]
  wire  _T_25; // @[LZD.scala 49:16]
  wire  _T_26; // @[LZD.scala 49:27]
  wire  _T_27; // @[LZD.scala 49:25]
  wire  _T_28; // @[LZD.scala 49:47]
  wire  _T_29; // @[LZD.scala 49:59]
  wire  _T_30; // @[LZD.scala 49:35]
  wire [2:0] _T_32; // @[Cat.scala 29:58]
  wire [3:0] _T_33; // @[LZD.scala 44:32]
  wire [1:0] _T_34; // @[LZD.scala 43:32]
  wire  _T_35; // @[LZD.scala 39:14]
  wire  _T_36; // @[LZD.scala 39:21]
  wire  _T_37; // @[LZD.scala 39:30]
  wire  _T_38; // @[LZD.scala 39:27]
  wire  _T_39; // @[LZD.scala 39:25]
  wire [1:0] _T_40; // @[Cat.scala 29:58]
  wire [1:0] _T_41; // @[LZD.scala 44:32]
  wire  _T_42; // @[LZD.scala 39:14]
  wire  _T_43; // @[LZD.scala 39:21]
  wire  _T_44; // @[LZD.scala 39:30]
  wire  _T_45; // @[LZD.scala 39:27]
  wire  _T_46; // @[LZD.scala 39:25]
  wire [1:0] _T_47; // @[Cat.scala 29:58]
  wire  _T_48; // @[Shift.scala 12:21]
  wire  _T_49; // @[Shift.scala 12:21]
  wire  _T_50; // @[LZD.scala 49:16]
  wire  _T_51; // @[LZD.scala 49:27]
  wire  _T_52; // @[LZD.scala 49:25]
  wire  _T_53; // @[LZD.scala 49:47]
  wire  _T_54; // @[LZD.scala 49:59]
  wire  _T_55; // @[LZD.scala 49:35]
  wire [2:0] _T_57; // @[Cat.scala 29:58]
  wire  _T_58; // @[Shift.scala 12:21]
  wire  _T_59; // @[Shift.scala 12:21]
  wire  _T_60; // @[LZD.scala 49:16]
  wire  _T_61; // @[LZD.scala 49:27]
  wire  _T_62; // @[LZD.scala 49:25]
  wire [1:0] _T_63; // @[LZD.scala 49:47]
  wire [1:0] _T_64; // @[LZD.scala 49:59]
  wire [1:0] _T_65; // @[LZD.scala 49:35]
  wire [3:0] _T_67; // @[Cat.scala 29:58]
  wire [5:0] _T_68; // @[LZD.scala 44:32]
  wire [3:0] _T_69; // @[LZD.scala 43:32]
  wire [1:0] _T_70; // @[LZD.scala 43:32]
  wire  _T_71; // @[LZD.scala 39:14]
  wire  _T_72; // @[LZD.scala 39:21]
  wire  _T_73; // @[LZD.scala 39:30]
  wire  _T_74; // @[LZD.scala 39:27]
  wire  _T_75; // @[LZD.scala 39:25]
  wire [1:0] _T_76; // @[Cat.scala 29:58]
  wire [1:0] _T_77; // @[LZD.scala 44:32]
  wire  _T_78; // @[LZD.scala 39:14]
  wire  _T_79; // @[LZD.scala 39:21]
  wire  _T_80; // @[LZD.scala 39:30]
  wire  _T_81; // @[LZD.scala 39:27]
  wire  _T_82; // @[LZD.scala 39:25]
  wire [1:0] _T_83; // @[Cat.scala 29:58]
  wire  _T_84; // @[Shift.scala 12:21]
  wire  _T_85; // @[Shift.scala 12:21]
  wire  _T_86; // @[LZD.scala 49:16]
  wire  _T_87; // @[LZD.scala 49:27]
  wire  _T_88; // @[LZD.scala 49:25]
  wire  _T_89; // @[LZD.scala 49:47]
  wire  _T_90; // @[LZD.scala 49:59]
  wire  _T_91; // @[LZD.scala 49:35]
  wire [2:0] _T_93; // @[Cat.scala 29:58]
  wire [1:0] _T_94; // @[LZD.scala 44:32]
  wire  _T_95; // @[LZD.scala 39:14]
  wire  _T_96; // @[LZD.scala 39:21]
  wire  _T_97; // @[LZD.scala 39:30]
  wire  _T_98; // @[LZD.scala 39:27]
  wire  _T_99; // @[LZD.scala 39:25]
  wire [1:0] _T_100; // @[Cat.scala 29:58]
  wire  _T_101; // @[Shift.scala 12:21]
  wire [1:0] _T_103; // @[LZD.scala 55:32]
  wire [1:0] _T_104; // @[LZD.scala 55:20]
  wire [2:0] _T_105; // @[Cat.scala 29:58]
  wire  _T_106; // @[Shift.scala 12:21]
  wire [2:0] _T_108; // @[LZD.scala 55:32]
  wire [2:0] _T_109; // @[LZD.scala 55:20]
  wire [3:0] _T_110; // @[Cat.scala 29:58]
  wire [3:0] _T_111; // @[convert.scala 21:22]
  wire [12:0] _T_112; // @[convert.scala 22:36]
  wire  _T_113; // @[Shift.scala 16:24]
  wire  _T_115; // @[Shift.scala 12:21]
  wire [4:0] _T_116; // @[Shift.scala 64:52]
  wire [12:0] _T_118; // @[Cat.scala 29:58]
  wire [12:0] _T_119; // @[Shift.scala 64:27]
  wire [2:0] _T_120; // @[Shift.scala 66:70]
  wire  _T_121; // @[Shift.scala 12:21]
  wire [8:0] _T_122; // @[Shift.scala 64:52]
  wire [12:0] _T_124; // @[Cat.scala 29:58]
  wire [12:0] _T_125; // @[Shift.scala 64:27]
  wire [1:0] _T_126; // @[Shift.scala 66:70]
  wire  _T_127; // @[Shift.scala 12:21]
  wire [10:0] _T_128; // @[Shift.scala 64:52]
  wire [12:0] _T_130; // @[Cat.scala 29:58]
  wire [12:0] _T_131; // @[Shift.scala 64:27]
  wire  _T_132; // @[Shift.scala 66:70]
  wire [11:0] _T_134; // @[Shift.scala 64:52]
  wire [12:0] _T_135; // @[Cat.scala 29:58]
  wire [12:0] _T_136; // @[Shift.scala 64:27]
  wire [12:0] _T_137; // @[Shift.scala 16:10]
  wire [2:0] _T_138; // @[convert.scala 23:34]
  wire [9:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_140; // @[convert.scala 25:26]
  wire [3:0] _T_142; // @[convert.scala 25:42]
  wire [2:0] _T_145; // @[convert.scala 26:67]
  wire [2:0] _T_146; // @[convert.scala 26:51]
  wire [7:0] _T_147; // @[Cat.scala 29:58]
  wire [14:0] _T_149; // @[convert.scala 29:56]
  wire  _T_150; // @[convert.scala 29:60]
  wire  _T_151; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_154; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [7:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_163; // @[convert.scala 18:24]
  wire  _T_164; // @[convert.scala 18:40]
  wire  _T_165; // @[convert.scala 18:36]
  wire [13:0] _T_166; // @[convert.scala 19:24]
  wire [13:0] _T_167; // @[convert.scala 19:43]
  wire [13:0] _T_168; // @[convert.scala 19:39]
  wire [7:0] _T_169; // @[LZD.scala 43:32]
  wire [3:0] _T_170; // @[LZD.scala 43:32]
  wire [1:0] _T_171; // @[LZD.scala 43:32]
  wire  _T_172; // @[LZD.scala 39:14]
  wire  _T_173; // @[LZD.scala 39:21]
  wire  _T_174; // @[LZD.scala 39:30]
  wire  _T_175; // @[LZD.scala 39:27]
  wire  _T_176; // @[LZD.scala 39:25]
  wire [1:0] _T_177; // @[Cat.scala 29:58]
  wire [1:0] _T_178; // @[LZD.scala 44:32]
  wire  _T_179; // @[LZD.scala 39:14]
  wire  _T_180; // @[LZD.scala 39:21]
  wire  _T_181; // @[LZD.scala 39:30]
  wire  _T_182; // @[LZD.scala 39:27]
  wire  _T_183; // @[LZD.scala 39:25]
  wire [1:0] _T_184; // @[Cat.scala 29:58]
  wire  _T_185; // @[Shift.scala 12:21]
  wire  _T_186; // @[Shift.scala 12:21]
  wire  _T_187; // @[LZD.scala 49:16]
  wire  _T_188; // @[LZD.scala 49:27]
  wire  _T_189; // @[LZD.scala 49:25]
  wire  _T_190; // @[LZD.scala 49:47]
  wire  _T_191; // @[LZD.scala 49:59]
  wire  _T_192; // @[LZD.scala 49:35]
  wire [2:0] _T_194; // @[Cat.scala 29:58]
  wire [3:0] _T_195; // @[LZD.scala 44:32]
  wire [1:0] _T_196; // @[LZD.scala 43:32]
  wire  _T_197; // @[LZD.scala 39:14]
  wire  _T_198; // @[LZD.scala 39:21]
  wire  _T_199; // @[LZD.scala 39:30]
  wire  _T_200; // @[LZD.scala 39:27]
  wire  _T_201; // @[LZD.scala 39:25]
  wire [1:0] _T_202; // @[Cat.scala 29:58]
  wire [1:0] _T_203; // @[LZD.scala 44:32]
  wire  _T_204; // @[LZD.scala 39:14]
  wire  _T_205; // @[LZD.scala 39:21]
  wire  _T_206; // @[LZD.scala 39:30]
  wire  _T_207; // @[LZD.scala 39:27]
  wire  _T_208; // @[LZD.scala 39:25]
  wire [1:0] _T_209; // @[Cat.scala 29:58]
  wire  _T_210; // @[Shift.scala 12:21]
  wire  _T_211; // @[Shift.scala 12:21]
  wire  _T_212; // @[LZD.scala 49:16]
  wire  _T_213; // @[LZD.scala 49:27]
  wire  _T_214; // @[LZD.scala 49:25]
  wire  _T_215; // @[LZD.scala 49:47]
  wire  _T_216; // @[LZD.scala 49:59]
  wire  _T_217; // @[LZD.scala 49:35]
  wire [2:0] _T_219; // @[Cat.scala 29:58]
  wire  _T_220; // @[Shift.scala 12:21]
  wire  _T_221; // @[Shift.scala 12:21]
  wire  _T_222; // @[LZD.scala 49:16]
  wire  _T_223; // @[LZD.scala 49:27]
  wire  _T_224; // @[LZD.scala 49:25]
  wire [1:0] _T_225; // @[LZD.scala 49:47]
  wire [1:0] _T_226; // @[LZD.scala 49:59]
  wire [1:0] _T_227; // @[LZD.scala 49:35]
  wire [3:0] _T_229; // @[Cat.scala 29:58]
  wire [5:0] _T_230; // @[LZD.scala 44:32]
  wire [3:0] _T_231; // @[LZD.scala 43:32]
  wire [1:0] _T_232; // @[LZD.scala 43:32]
  wire  _T_233; // @[LZD.scala 39:14]
  wire  _T_234; // @[LZD.scala 39:21]
  wire  _T_235; // @[LZD.scala 39:30]
  wire  _T_236; // @[LZD.scala 39:27]
  wire  _T_237; // @[LZD.scala 39:25]
  wire [1:0] _T_238; // @[Cat.scala 29:58]
  wire [1:0] _T_239; // @[LZD.scala 44:32]
  wire  _T_240; // @[LZD.scala 39:14]
  wire  _T_241; // @[LZD.scala 39:21]
  wire  _T_242; // @[LZD.scala 39:30]
  wire  _T_243; // @[LZD.scala 39:27]
  wire  _T_244; // @[LZD.scala 39:25]
  wire [1:0] _T_245; // @[Cat.scala 29:58]
  wire  _T_246; // @[Shift.scala 12:21]
  wire  _T_247; // @[Shift.scala 12:21]
  wire  _T_248; // @[LZD.scala 49:16]
  wire  _T_249; // @[LZD.scala 49:27]
  wire  _T_250; // @[LZD.scala 49:25]
  wire  _T_251; // @[LZD.scala 49:47]
  wire  _T_252; // @[LZD.scala 49:59]
  wire  _T_253; // @[LZD.scala 49:35]
  wire [2:0] _T_255; // @[Cat.scala 29:58]
  wire [1:0] _T_256; // @[LZD.scala 44:32]
  wire  _T_257; // @[LZD.scala 39:14]
  wire  _T_258; // @[LZD.scala 39:21]
  wire  _T_259; // @[LZD.scala 39:30]
  wire  _T_260; // @[LZD.scala 39:27]
  wire  _T_261; // @[LZD.scala 39:25]
  wire [1:0] _T_262; // @[Cat.scala 29:58]
  wire  _T_263; // @[Shift.scala 12:21]
  wire [1:0] _T_265; // @[LZD.scala 55:32]
  wire [1:0] _T_266; // @[LZD.scala 55:20]
  wire [2:0] _T_267; // @[Cat.scala 29:58]
  wire  _T_268; // @[Shift.scala 12:21]
  wire [2:0] _T_270; // @[LZD.scala 55:32]
  wire [2:0] _T_271; // @[LZD.scala 55:20]
  wire [3:0] _T_272; // @[Cat.scala 29:58]
  wire [3:0] _T_273; // @[convert.scala 21:22]
  wire [12:0] _T_274; // @[convert.scala 22:36]
  wire  _T_275; // @[Shift.scala 16:24]
  wire  _T_277; // @[Shift.scala 12:21]
  wire [4:0] _T_278; // @[Shift.scala 64:52]
  wire [12:0] _T_280; // @[Cat.scala 29:58]
  wire [12:0] _T_281; // @[Shift.scala 64:27]
  wire [2:0] _T_282; // @[Shift.scala 66:70]
  wire  _T_283; // @[Shift.scala 12:21]
  wire [8:0] _T_284; // @[Shift.scala 64:52]
  wire [12:0] _T_286; // @[Cat.scala 29:58]
  wire [12:0] _T_287; // @[Shift.scala 64:27]
  wire [1:0] _T_288; // @[Shift.scala 66:70]
  wire  _T_289; // @[Shift.scala 12:21]
  wire [10:0] _T_290; // @[Shift.scala 64:52]
  wire [12:0] _T_292; // @[Cat.scala 29:58]
  wire [12:0] _T_293; // @[Shift.scala 64:27]
  wire  _T_294; // @[Shift.scala 66:70]
  wire [11:0] _T_296; // @[Shift.scala 64:52]
  wire [12:0] _T_297; // @[Cat.scala 29:58]
  wire [12:0] _T_298; // @[Shift.scala 64:27]
  wire [12:0] _T_299; // @[Shift.scala 16:10]
  wire [2:0] _T_300; // @[convert.scala 23:34]
  wire [9:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_302; // @[convert.scala 25:26]
  wire [3:0] _T_304; // @[convert.scala 25:42]
  wire [2:0] _T_307; // @[convert.scala 26:67]
  wire [2:0] _T_308; // @[convert.scala 26:51]
  wire [7:0] _T_309; // @[Cat.scala 29:58]
  wire [14:0] _T_311; // @[convert.scala 29:56]
  wire  _T_312; // @[convert.scala 29:60]
  wire  _T_313; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_316; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [7:0] decB_scale; // @[convert.scala 32:24]
  wire  aGTb; // @[PositAdder.scala 24:32]
  wire  greaterSign; // @[PositAdder.scala 25:24]
  wire  smallerSign; // @[PositAdder.scala 26:24]
  wire [7:0] greaterExp; // @[PositAdder.scala 27:24]
  wire [7:0] smallerExp; // @[PositAdder.scala 28:24]
  wire [9:0] greaterFrac; // @[PositAdder.scala 29:24]
  wire [9:0] smallerFrac; // @[PositAdder.scala 30:24]
  wire  smallerZero; // @[PositAdder.scala 31:24]
  wire [7:0] _T_325; // @[PositAdder.scala 32:32]
  wire [7:0] scale_diff; // @[PositAdder.scala 32:32]
  wire  _T_326; // @[PositAdder.scala 33:38]
  wire [11:0] greaterSig; // @[Cat.scala 29:58]
  wire  _T_328; // @[PositAdder.scala 34:52]
  wire  _T_329; // @[PositAdder.scala 34:38]
  wire [14:0] _T_332; // @[Cat.scala 29:58]
  wire [7:0] _T_333; // @[PositAdder.scala 35:68]
  wire  _T_334; // @[Shift.scala 39:24]
  wire [3:0] _T_335; // @[Shift.scala 40:44]
  wire [6:0] _T_336; // @[Shift.scala 90:30]
  wire [7:0] _T_337; // @[Shift.scala 90:48]
  wire  _T_338; // @[Shift.scala 90:57]
  wire [6:0] _GEN_0; // @[Shift.scala 90:39]
  wire [6:0] _T_339; // @[Shift.scala 90:39]
  wire  _T_340; // @[Shift.scala 12:21]
  wire  _T_341; // @[Shift.scala 12:21]
  wire [7:0] _T_343; // @[Bitwise.scala 71:12]
  wire [14:0] _T_344; // @[Cat.scala 29:58]
  wire [14:0] _T_345; // @[Shift.scala 91:22]
  wire [2:0] _T_346; // @[Shift.scala 92:77]
  wire [10:0] _T_347; // @[Shift.scala 90:30]
  wire [3:0] _T_348; // @[Shift.scala 90:48]
  wire  _T_349; // @[Shift.scala 90:57]
  wire [10:0] _GEN_1; // @[Shift.scala 90:39]
  wire [10:0] _T_350; // @[Shift.scala 90:39]
  wire  _T_351; // @[Shift.scala 12:21]
  wire  _T_352; // @[Shift.scala 12:21]
  wire [3:0] _T_354; // @[Bitwise.scala 71:12]
  wire [14:0] _T_355; // @[Cat.scala 29:58]
  wire [14:0] _T_356; // @[Shift.scala 91:22]
  wire [1:0] _T_357; // @[Shift.scala 92:77]
  wire [12:0] _T_358; // @[Shift.scala 90:30]
  wire [1:0] _T_359; // @[Shift.scala 90:48]
  wire  _T_360; // @[Shift.scala 90:57]
  wire [12:0] _GEN_2; // @[Shift.scala 90:39]
  wire [12:0] _T_361; // @[Shift.scala 90:39]
  wire  _T_362; // @[Shift.scala 12:21]
  wire  _T_363; // @[Shift.scala 12:21]
  wire [1:0] _T_365; // @[Bitwise.scala 71:12]
  wire [14:0] _T_366; // @[Cat.scala 29:58]
  wire [14:0] _T_367; // @[Shift.scala 91:22]
  wire  _T_368; // @[Shift.scala 92:77]
  wire [13:0] _T_369; // @[Shift.scala 90:30]
  wire  _T_370; // @[Shift.scala 90:48]
  wire [13:0] _GEN_3; // @[Shift.scala 90:39]
  wire [13:0] _T_372; // @[Shift.scala 90:39]
  wire  _T_374; // @[Shift.scala 12:21]
  wire [14:0] _T_375; // @[Cat.scala 29:58]
  wire [14:0] _T_376; // @[Shift.scala 91:22]
  wire [14:0] _T_379; // @[Bitwise.scala 71:12]
  wire [14:0] smallerSig; // @[Shift.scala 39:10]
  wire [11:0] _T_380; // @[PositAdder.scala 36:45]
  wire [12:0] rawSumSig; // @[PositAdder.scala 36:32]
  wire  _T_381; // @[PositAdder.scala 37:31]
  wire  _T_382; // @[PositAdder.scala 37:59]
  wire  sumSign; // @[PositAdder.scala 37:43]
  wire [11:0] _T_383; // @[PositAdder.scala 38:48]
  wire [2:0] _T_384; // @[PositAdder.scala 38:63]
  wire [15:0] signSumSig; // @[Cat.scala 29:58]
  wire [14:0] _T_386; // @[PositAdder.scala 40:31]
  wire [14:0] _T_387; // @[PositAdder.scala 40:66]
  wire [14:0] sumXor; // @[PositAdder.scala 40:49]
  wire [7:0] _T_388; // @[LZD.scala 43:32]
  wire [3:0] _T_389; // @[LZD.scala 43:32]
  wire [1:0] _T_390; // @[LZD.scala 43:32]
  wire  _T_391; // @[LZD.scala 39:14]
  wire  _T_392; // @[LZD.scala 39:21]
  wire  _T_393; // @[LZD.scala 39:30]
  wire  _T_394; // @[LZD.scala 39:27]
  wire  _T_395; // @[LZD.scala 39:25]
  wire [1:0] _T_396; // @[Cat.scala 29:58]
  wire [1:0] _T_397; // @[LZD.scala 44:32]
  wire  _T_398; // @[LZD.scala 39:14]
  wire  _T_399; // @[LZD.scala 39:21]
  wire  _T_400; // @[LZD.scala 39:30]
  wire  _T_401; // @[LZD.scala 39:27]
  wire  _T_402; // @[LZD.scala 39:25]
  wire [1:0] _T_403; // @[Cat.scala 29:58]
  wire  _T_404; // @[Shift.scala 12:21]
  wire  _T_405; // @[Shift.scala 12:21]
  wire  _T_406; // @[LZD.scala 49:16]
  wire  _T_407; // @[LZD.scala 49:27]
  wire  _T_408; // @[LZD.scala 49:25]
  wire  _T_409; // @[LZD.scala 49:47]
  wire  _T_410; // @[LZD.scala 49:59]
  wire  _T_411; // @[LZD.scala 49:35]
  wire [2:0] _T_413; // @[Cat.scala 29:58]
  wire [3:0] _T_414; // @[LZD.scala 44:32]
  wire [1:0] _T_415; // @[LZD.scala 43:32]
  wire  _T_416; // @[LZD.scala 39:14]
  wire  _T_417; // @[LZD.scala 39:21]
  wire  _T_418; // @[LZD.scala 39:30]
  wire  _T_419; // @[LZD.scala 39:27]
  wire  _T_420; // @[LZD.scala 39:25]
  wire [1:0] _T_421; // @[Cat.scala 29:58]
  wire [1:0] _T_422; // @[LZD.scala 44:32]
  wire  _T_423; // @[LZD.scala 39:14]
  wire  _T_424; // @[LZD.scala 39:21]
  wire  _T_425; // @[LZD.scala 39:30]
  wire  _T_426; // @[LZD.scala 39:27]
  wire  _T_427; // @[LZD.scala 39:25]
  wire [1:0] _T_428; // @[Cat.scala 29:58]
  wire  _T_429; // @[Shift.scala 12:21]
  wire  _T_430; // @[Shift.scala 12:21]
  wire  _T_431; // @[LZD.scala 49:16]
  wire  _T_432; // @[LZD.scala 49:27]
  wire  _T_433; // @[LZD.scala 49:25]
  wire  _T_434; // @[LZD.scala 49:47]
  wire  _T_435; // @[LZD.scala 49:59]
  wire  _T_436; // @[LZD.scala 49:35]
  wire [2:0] _T_438; // @[Cat.scala 29:58]
  wire  _T_439; // @[Shift.scala 12:21]
  wire  _T_440; // @[Shift.scala 12:21]
  wire  _T_441; // @[LZD.scala 49:16]
  wire  _T_442; // @[LZD.scala 49:27]
  wire  _T_443; // @[LZD.scala 49:25]
  wire [1:0] _T_444; // @[LZD.scala 49:47]
  wire [1:0] _T_445; // @[LZD.scala 49:59]
  wire [1:0] _T_446; // @[LZD.scala 49:35]
  wire [3:0] _T_448; // @[Cat.scala 29:58]
  wire [6:0] _T_449; // @[LZD.scala 44:32]
  wire [3:0] _T_450; // @[LZD.scala 43:32]
  wire [1:0] _T_451; // @[LZD.scala 43:32]
  wire  _T_452; // @[LZD.scala 39:14]
  wire  _T_453; // @[LZD.scala 39:21]
  wire  _T_454; // @[LZD.scala 39:30]
  wire  _T_455; // @[LZD.scala 39:27]
  wire  _T_456; // @[LZD.scala 39:25]
  wire [1:0] _T_457; // @[Cat.scala 29:58]
  wire [1:0] _T_458; // @[LZD.scala 44:32]
  wire  _T_459; // @[LZD.scala 39:14]
  wire  _T_460; // @[LZD.scala 39:21]
  wire  _T_461; // @[LZD.scala 39:30]
  wire  _T_462; // @[LZD.scala 39:27]
  wire  _T_463; // @[LZD.scala 39:25]
  wire [1:0] _T_464; // @[Cat.scala 29:58]
  wire  _T_465; // @[Shift.scala 12:21]
  wire  _T_466; // @[Shift.scala 12:21]
  wire  _T_467; // @[LZD.scala 49:16]
  wire  _T_468; // @[LZD.scala 49:27]
  wire  _T_469; // @[LZD.scala 49:25]
  wire  _T_470; // @[LZD.scala 49:47]
  wire  _T_471; // @[LZD.scala 49:59]
  wire  _T_472; // @[LZD.scala 49:35]
  wire [2:0] _T_474; // @[Cat.scala 29:58]
  wire [2:0] _T_475; // @[LZD.scala 44:32]
  wire [1:0] _T_476; // @[LZD.scala 43:32]
  wire  _T_477; // @[LZD.scala 39:14]
  wire  _T_478; // @[LZD.scala 39:21]
  wire  _T_479; // @[LZD.scala 39:30]
  wire  _T_480; // @[LZD.scala 39:27]
  wire  _T_481; // @[LZD.scala 39:25]
  wire [1:0] _T_482; // @[Cat.scala 29:58]
  wire  _T_483; // @[LZD.scala 44:32]
  wire  _T_485; // @[Shift.scala 12:21]
  wire  _T_487; // @[LZD.scala 55:32]
  wire  _T_488; // @[LZD.scala 55:20]
  wire [1:0] _T_489; // @[Cat.scala 29:58]
  wire  _T_490; // @[Shift.scala 12:21]
  wire [1:0] _T_492; // @[LZD.scala 55:32]
  wire [1:0] _T_493; // @[LZD.scala 55:20]
  wire [2:0] _T_494; // @[Cat.scala 29:58]
  wire  _T_495; // @[Shift.scala 12:21]
  wire [2:0] _T_497; // @[LZD.scala 55:32]
  wire [2:0] _T_498; // @[LZD.scala 55:20]
  wire [3:0] sumLZD; // @[Cat.scala 29:58]
  wire [4:0] _T_499; // @[Cat.scala 29:58]
  wire [4:0] _T_500; // @[PositAdder.scala 42:38]
  wire [4:0] _T_502; // @[PositAdder.scala 42:45]
  wire [4:0] scaleBias; // @[PositAdder.scala 42:45]
  wire [7:0] _GEN_4; // @[PositAdder.scala 43:32]
  wire [8:0] sumScale; // @[PositAdder.scala 43:32]
  wire  overflow; // @[PositAdder.scala 44:30]
  wire [3:0] normalShift; // @[PositAdder.scala 45:22]
  wire [13:0] _T_503; // @[PositAdder.scala 46:36]
  wire  _T_504; // @[Shift.scala 16:24]
  wire  _T_506; // @[Shift.scala 12:21]
  wire [5:0] _T_507; // @[Shift.scala 64:52]
  wire [13:0] _T_509; // @[Cat.scala 29:58]
  wire [13:0] _T_510; // @[Shift.scala 64:27]
  wire [2:0] _T_511; // @[Shift.scala 66:70]
  wire  _T_512; // @[Shift.scala 12:21]
  wire [9:0] _T_513; // @[Shift.scala 64:52]
  wire [13:0] _T_515; // @[Cat.scala 29:58]
  wire [13:0] _T_516; // @[Shift.scala 64:27]
  wire [1:0] _T_517; // @[Shift.scala 66:70]
  wire  _T_518; // @[Shift.scala 12:21]
  wire [11:0] _T_519; // @[Shift.scala 64:52]
  wire [13:0] _T_521; // @[Cat.scala 29:58]
  wire [13:0] _T_522; // @[Shift.scala 64:27]
  wire  _T_523; // @[Shift.scala 66:70]
  wire [12:0] _T_525; // @[Shift.scala 64:52]
  wire [13:0] _T_526; // @[Cat.scala 29:58]
  wire [13:0] _T_527; // @[Shift.scala 64:27]
  wire [13:0] shiftSig; // @[Shift.scala 16:10]
  wire [8:0] _T_528; // @[PositAdder.scala 51:24]
  wire [9:0] decS_fraction; // @[PositAdder.scala 52:34]
  wire  decS_isNaR; // @[PositAdder.scala 53:32]
  wire  _T_531; // @[PositAdder.scala 54:33]
  wire  _T_532; // @[PositAdder.scala 54:21]
  wire  _T_533; // @[PositAdder.scala 54:52]
  wire  decS_isZero; // @[PositAdder.scala 54:37]
  wire [1:0] _T_535; // @[PositAdder.scala 55:33]
  wire  _T_536; // @[PositAdder.scala 55:49]
  wire  _T_537; // @[PositAdder.scala 55:63]
  wire  _T_538; // @[PositAdder.scala 55:53]
  wire [7:0] _GEN_5; // @[PositAdder.scala 48:25 PositAdder.scala 51:18]
  wire [7:0] decS_scale; // @[PositAdder.scala 48:25 PositAdder.scala 51:18]
  wire [2:0] _T_541; // @[convert.scala 46:61]
  wire [2:0] _T_542; // @[convert.scala 46:52]
  wire [2:0] _T_544; // @[convert.scala 46:42]
  wire [4:0] _T_545; // @[convert.scala 48:34]
  wire  _T_546; // @[convert.scala 49:36]
  wire [4:0] _T_548; // @[convert.scala 50:36]
  wire [4:0] _T_549; // @[convert.scala 50:36]
  wire [4:0] _T_550; // @[convert.scala 50:28]
  wire  _T_551; // @[convert.scala 51:31]
  wire  _T_552; // @[convert.scala 52:43]
  wire [17:0] _T_556; // @[Cat.scala 29:58]
  wire [4:0] _T_557; // @[Shift.scala 39:17]
  wire  _T_558; // @[Shift.scala 39:24]
  wire [1:0] _T_560; // @[Shift.scala 90:30]
  wire [15:0] _T_561; // @[Shift.scala 90:48]
  wire  _T_562; // @[Shift.scala 90:57]
  wire [1:0] _GEN_6; // @[Shift.scala 90:39]
  wire [1:0] _T_563; // @[Shift.scala 90:39]
  wire  _T_564; // @[Shift.scala 12:21]
  wire  _T_565; // @[Shift.scala 12:21]
  wire [15:0] _T_567; // @[Bitwise.scala 71:12]
  wire [17:0] _T_568; // @[Cat.scala 29:58]
  wire [17:0] _T_569; // @[Shift.scala 91:22]
  wire [3:0] _T_570; // @[Shift.scala 92:77]
  wire [9:0] _T_571; // @[Shift.scala 90:30]
  wire [7:0] _T_572; // @[Shift.scala 90:48]
  wire  _T_573; // @[Shift.scala 90:57]
  wire [9:0] _GEN_7; // @[Shift.scala 90:39]
  wire [9:0] _T_574; // @[Shift.scala 90:39]
  wire  _T_575; // @[Shift.scala 12:21]
  wire  _T_576; // @[Shift.scala 12:21]
  wire [7:0] _T_578; // @[Bitwise.scala 71:12]
  wire [17:0] _T_579; // @[Cat.scala 29:58]
  wire [17:0] _T_580; // @[Shift.scala 91:22]
  wire [2:0] _T_581; // @[Shift.scala 92:77]
  wire [13:0] _T_582; // @[Shift.scala 90:30]
  wire [3:0] _T_583; // @[Shift.scala 90:48]
  wire  _T_584; // @[Shift.scala 90:57]
  wire [13:0] _GEN_8; // @[Shift.scala 90:39]
  wire [13:0] _T_585; // @[Shift.scala 90:39]
  wire  _T_586; // @[Shift.scala 12:21]
  wire  _T_587; // @[Shift.scala 12:21]
  wire [3:0] _T_589; // @[Bitwise.scala 71:12]
  wire [17:0] _T_590; // @[Cat.scala 29:58]
  wire [17:0] _T_591; // @[Shift.scala 91:22]
  wire [1:0] _T_592; // @[Shift.scala 92:77]
  wire [15:0] _T_593; // @[Shift.scala 90:30]
  wire [1:0] _T_594; // @[Shift.scala 90:48]
  wire  _T_595; // @[Shift.scala 90:57]
  wire [15:0] _GEN_9; // @[Shift.scala 90:39]
  wire [15:0] _T_596; // @[Shift.scala 90:39]
  wire  _T_597; // @[Shift.scala 12:21]
  wire  _T_598; // @[Shift.scala 12:21]
  wire [1:0] _T_600; // @[Bitwise.scala 71:12]
  wire [17:0] _T_601; // @[Cat.scala 29:58]
  wire [17:0] _T_602; // @[Shift.scala 91:22]
  wire  _T_603; // @[Shift.scala 92:77]
  wire [16:0] _T_604; // @[Shift.scala 90:30]
  wire  _T_605; // @[Shift.scala 90:48]
  wire [16:0] _GEN_10; // @[Shift.scala 90:39]
  wire [16:0] _T_607; // @[Shift.scala 90:39]
  wire  _T_609; // @[Shift.scala 12:21]
  wire [17:0] _T_610; // @[Cat.scala 29:58]
  wire [17:0] _T_611; // @[Shift.scala 91:22]
  wire [17:0] _T_614; // @[Bitwise.scala 71:12]
  wire [17:0] _T_615; // @[Shift.scala 39:10]
  wire  _T_616; // @[convert.scala 55:31]
  wire  _T_617; // @[convert.scala 56:31]
  wire  _T_618; // @[convert.scala 57:31]
  wire  _T_619; // @[convert.scala 58:31]
  wire [14:0] _T_620; // @[convert.scala 59:69]
  wire  _T_621; // @[convert.scala 59:81]
  wire  _T_622; // @[convert.scala 59:50]
  wire  _T_624; // @[convert.scala 60:81]
  wire  _T_625; // @[convert.scala 61:44]
  wire  _T_626; // @[convert.scala 61:52]
  wire  _T_627; // @[convert.scala 61:36]
  wire  _T_628; // @[convert.scala 62:63]
  wire  _T_629; // @[convert.scala 62:103]
  wire  _T_630; // @[convert.scala 62:60]
  wire [14:0] _GEN_11; // @[convert.scala 63:56]
  wire [14:0] _T_633; // @[convert.scala 63:56]
  wire [15:0] _T_634; // @[Cat.scala 29:58]
  wire [15:0] _T_636; // @[Mux.scala 87:16]
  assign _T_1 = io_A[15]; // @[convert.scala 18:24]
  assign _T_2 = io_A[14]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[14:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[13:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[13:6]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[7:4]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8[3:2]; // @[LZD.scala 43:32]
  assign _T_10 = _T_9 != 2'h0; // @[LZD.scala 39:14]
  assign _T_11 = _T_9[1]; // @[LZD.scala 39:21]
  assign _T_12 = _T_9[0]; // @[LZD.scala 39:30]
  assign _T_13 = ~ _T_12; // @[LZD.scala 39:27]
  assign _T_14 = _T_11 | _T_13; // @[LZD.scala 39:25]
  assign _T_15 = {_T_10,_T_14}; // @[Cat.scala 29:58]
  assign _T_16 = _T_8[1:0]; // @[LZD.scala 44:32]
  assign _T_17 = _T_16 != 2'h0; // @[LZD.scala 39:14]
  assign _T_18 = _T_16[1]; // @[LZD.scala 39:21]
  assign _T_19 = _T_16[0]; // @[LZD.scala 39:30]
  assign _T_20 = ~ _T_19; // @[LZD.scala 39:27]
  assign _T_21 = _T_18 | _T_20; // @[LZD.scala 39:25]
  assign _T_22 = {_T_17,_T_21}; // @[Cat.scala 29:58]
  assign _T_23 = _T_15[1]; // @[Shift.scala 12:21]
  assign _T_24 = _T_22[1]; // @[Shift.scala 12:21]
  assign _T_25 = _T_23 | _T_24; // @[LZD.scala 49:16]
  assign _T_26 = ~ _T_24; // @[LZD.scala 49:27]
  assign _T_27 = _T_23 | _T_26; // @[LZD.scala 49:25]
  assign _T_28 = _T_15[0:0]; // @[LZD.scala 49:47]
  assign _T_29 = _T_22[0:0]; // @[LZD.scala 49:59]
  assign _T_30 = _T_23 ? _T_28 : _T_29; // @[LZD.scala 49:35]
  assign _T_32 = {_T_25,_T_27,_T_30}; // @[Cat.scala 29:58]
  assign _T_33 = _T_7[3:0]; // @[LZD.scala 44:32]
  assign _T_34 = _T_33[3:2]; // @[LZD.scala 43:32]
  assign _T_35 = _T_34 != 2'h0; // @[LZD.scala 39:14]
  assign _T_36 = _T_34[1]; // @[LZD.scala 39:21]
  assign _T_37 = _T_34[0]; // @[LZD.scala 39:30]
  assign _T_38 = ~ _T_37; // @[LZD.scala 39:27]
  assign _T_39 = _T_36 | _T_38; // @[LZD.scala 39:25]
  assign _T_40 = {_T_35,_T_39}; // @[Cat.scala 29:58]
  assign _T_41 = _T_33[1:0]; // @[LZD.scala 44:32]
  assign _T_42 = _T_41 != 2'h0; // @[LZD.scala 39:14]
  assign _T_43 = _T_41[1]; // @[LZD.scala 39:21]
  assign _T_44 = _T_41[0]; // @[LZD.scala 39:30]
  assign _T_45 = ~ _T_44; // @[LZD.scala 39:27]
  assign _T_46 = _T_43 | _T_45; // @[LZD.scala 39:25]
  assign _T_47 = {_T_42,_T_46}; // @[Cat.scala 29:58]
  assign _T_48 = _T_40[1]; // @[Shift.scala 12:21]
  assign _T_49 = _T_47[1]; // @[Shift.scala 12:21]
  assign _T_50 = _T_48 | _T_49; // @[LZD.scala 49:16]
  assign _T_51 = ~ _T_49; // @[LZD.scala 49:27]
  assign _T_52 = _T_48 | _T_51; // @[LZD.scala 49:25]
  assign _T_53 = _T_40[0:0]; // @[LZD.scala 49:47]
  assign _T_54 = _T_47[0:0]; // @[LZD.scala 49:59]
  assign _T_55 = _T_48 ? _T_53 : _T_54; // @[LZD.scala 49:35]
  assign _T_57 = {_T_50,_T_52,_T_55}; // @[Cat.scala 29:58]
  assign _T_58 = _T_32[2]; // @[Shift.scala 12:21]
  assign _T_59 = _T_57[2]; // @[Shift.scala 12:21]
  assign _T_60 = _T_58 | _T_59; // @[LZD.scala 49:16]
  assign _T_61 = ~ _T_59; // @[LZD.scala 49:27]
  assign _T_62 = _T_58 | _T_61; // @[LZD.scala 49:25]
  assign _T_63 = _T_32[1:0]; // @[LZD.scala 49:47]
  assign _T_64 = _T_57[1:0]; // @[LZD.scala 49:59]
  assign _T_65 = _T_58 ? _T_63 : _T_64; // @[LZD.scala 49:35]
  assign _T_67 = {_T_60,_T_62,_T_65}; // @[Cat.scala 29:58]
  assign _T_68 = _T_6[5:0]; // @[LZD.scala 44:32]
  assign _T_69 = _T_68[5:2]; // @[LZD.scala 43:32]
  assign _T_70 = _T_69[3:2]; // @[LZD.scala 43:32]
  assign _T_71 = _T_70 != 2'h0; // @[LZD.scala 39:14]
  assign _T_72 = _T_70[1]; // @[LZD.scala 39:21]
  assign _T_73 = _T_70[0]; // @[LZD.scala 39:30]
  assign _T_74 = ~ _T_73; // @[LZD.scala 39:27]
  assign _T_75 = _T_72 | _T_74; // @[LZD.scala 39:25]
  assign _T_76 = {_T_71,_T_75}; // @[Cat.scala 29:58]
  assign _T_77 = _T_69[1:0]; // @[LZD.scala 44:32]
  assign _T_78 = _T_77 != 2'h0; // @[LZD.scala 39:14]
  assign _T_79 = _T_77[1]; // @[LZD.scala 39:21]
  assign _T_80 = _T_77[0]; // @[LZD.scala 39:30]
  assign _T_81 = ~ _T_80; // @[LZD.scala 39:27]
  assign _T_82 = _T_79 | _T_81; // @[LZD.scala 39:25]
  assign _T_83 = {_T_78,_T_82}; // @[Cat.scala 29:58]
  assign _T_84 = _T_76[1]; // @[Shift.scala 12:21]
  assign _T_85 = _T_83[1]; // @[Shift.scala 12:21]
  assign _T_86 = _T_84 | _T_85; // @[LZD.scala 49:16]
  assign _T_87 = ~ _T_85; // @[LZD.scala 49:27]
  assign _T_88 = _T_84 | _T_87; // @[LZD.scala 49:25]
  assign _T_89 = _T_76[0:0]; // @[LZD.scala 49:47]
  assign _T_90 = _T_83[0:0]; // @[LZD.scala 49:59]
  assign _T_91 = _T_84 ? _T_89 : _T_90; // @[LZD.scala 49:35]
  assign _T_93 = {_T_86,_T_88,_T_91}; // @[Cat.scala 29:58]
  assign _T_94 = _T_68[1:0]; // @[LZD.scala 44:32]
  assign _T_95 = _T_94 != 2'h0; // @[LZD.scala 39:14]
  assign _T_96 = _T_94[1]; // @[LZD.scala 39:21]
  assign _T_97 = _T_94[0]; // @[LZD.scala 39:30]
  assign _T_98 = ~ _T_97; // @[LZD.scala 39:27]
  assign _T_99 = _T_96 | _T_98; // @[LZD.scala 39:25]
  assign _T_100 = {_T_95,_T_99}; // @[Cat.scala 29:58]
  assign _T_101 = _T_93[2]; // @[Shift.scala 12:21]
  assign _T_103 = _T_93[1:0]; // @[LZD.scala 55:32]
  assign _T_104 = _T_101 ? _T_103 : _T_100; // @[LZD.scala 55:20]
  assign _T_105 = {_T_101,_T_104}; // @[Cat.scala 29:58]
  assign _T_106 = _T_67[3]; // @[Shift.scala 12:21]
  assign _T_108 = _T_67[2:0]; // @[LZD.scala 55:32]
  assign _T_109 = _T_106 ? _T_108 : _T_105; // @[LZD.scala 55:20]
  assign _T_110 = {_T_106,_T_109}; // @[Cat.scala 29:58]
  assign _T_111 = ~ _T_110; // @[convert.scala 21:22]
  assign _T_112 = io_A[12:0]; // @[convert.scala 22:36]
  assign _T_113 = _T_111 < 4'hd; // @[Shift.scala 16:24]
  assign _T_115 = _T_111[3]; // @[Shift.scala 12:21]
  assign _T_116 = _T_112[4:0]; // @[Shift.scala 64:52]
  assign _T_118 = {_T_116,8'h0}; // @[Cat.scala 29:58]
  assign _T_119 = _T_115 ? _T_118 : _T_112; // @[Shift.scala 64:27]
  assign _T_120 = _T_111[2:0]; // @[Shift.scala 66:70]
  assign _T_121 = _T_120[2]; // @[Shift.scala 12:21]
  assign _T_122 = _T_119[8:0]; // @[Shift.scala 64:52]
  assign _T_124 = {_T_122,4'h0}; // @[Cat.scala 29:58]
  assign _T_125 = _T_121 ? _T_124 : _T_119; // @[Shift.scala 64:27]
  assign _T_126 = _T_120[1:0]; // @[Shift.scala 66:70]
  assign _T_127 = _T_126[1]; // @[Shift.scala 12:21]
  assign _T_128 = _T_125[10:0]; // @[Shift.scala 64:52]
  assign _T_130 = {_T_128,2'h0}; // @[Cat.scala 29:58]
  assign _T_131 = _T_127 ? _T_130 : _T_125; // @[Shift.scala 64:27]
  assign _T_132 = _T_126[0:0]; // @[Shift.scala 66:70]
  assign _T_134 = _T_131[11:0]; // @[Shift.scala 64:52]
  assign _T_135 = {_T_134,1'h0}; // @[Cat.scala 29:58]
  assign _T_136 = _T_132 ? _T_135 : _T_131; // @[Shift.scala 64:27]
  assign _T_137 = _T_113 ? _T_136 : 13'h0; // @[Shift.scala 16:10]
  assign _T_138 = _T_137[12:10]; // @[convert.scala 23:34]
  assign decA_fraction = _T_137[9:0]; // @[convert.scala 24:34]
  assign _T_140 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_142 = _T_3 ? _T_111 : _T_110; // @[convert.scala 25:42]
  assign _T_145 = ~ _T_138; // @[convert.scala 26:67]
  assign _T_146 = _T_1 ? _T_145 : _T_138; // @[convert.scala 26:51]
  assign _T_147 = {_T_140,_T_142,_T_146}; // @[Cat.scala 29:58]
  assign _T_149 = io_A[14:0]; // @[convert.scala 29:56]
  assign _T_150 = _T_149 != 15'h0; // @[convert.scala 29:60]
  assign _T_151 = ~ _T_150; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_151; // @[convert.scala 29:39]
  assign _T_154 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_154 & _T_151; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_147); // @[convert.scala 32:24]
  assign _T_163 = io_B[15]; // @[convert.scala 18:24]
  assign _T_164 = io_B[14]; // @[convert.scala 18:40]
  assign _T_165 = _T_163 ^ _T_164; // @[convert.scala 18:36]
  assign _T_166 = io_B[14:1]; // @[convert.scala 19:24]
  assign _T_167 = io_B[13:0]; // @[convert.scala 19:43]
  assign _T_168 = _T_166 ^ _T_167; // @[convert.scala 19:39]
  assign _T_169 = _T_168[13:6]; // @[LZD.scala 43:32]
  assign _T_170 = _T_169[7:4]; // @[LZD.scala 43:32]
  assign _T_171 = _T_170[3:2]; // @[LZD.scala 43:32]
  assign _T_172 = _T_171 != 2'h0; // @[LZD.scala 39:14]
  assign _T_173 = _T_171[1]; // @[LZD.scala 39:21]
  assign _T_174 = _T_171[0]; // @[LZD.scala 39:30]
  assign _T_175 = ~ _T_174; // @[LZD.scala 39:27]
  assign _T_176 = _T_173 | _T_175; // @[LZD.scala 39:25]
  assign _T_177 = {_T_172,_T_176}; // @[Cat.scala 29:58]
  assign _T_178 = _T_170[1:0]; // @[LZD.scala 44:32]
  assign _T_179 = _T_178 != 2'h0; // @[LZD.scala 39:14]
  assign _T_180 = _T_178[1]; // @[LZD.scala 39:21]
  assign _T_181 = _T_178[0]; // @[LZD.scala 39:30]
  assign _T_182 = ~ _T_181; // @[LZD.scala 39:27]
  assign _T_183 = _T_180 | _T_182; // @[LZD.scala 39:25]
  assign _T_184 = {_T_179,_T_183}; // @[Cat.scala 29:58]
  assign _T_185 = _T_177[1]; // @[Shift.scala 12:21]
  assign _T_186 = _T_184[1]; // @[Shift.scala 12:21]
  assign _T_187 = _T_185 | _T_186; // @[LZD.scala 49:16]
  assign _T_188 = ~ _T_186; // @[LZD.scala 49:27]
  assign _T_189 = _T_185 | _T_188; // @[LZD.scala 49:25]
  assign _T_190 = _T_177[0:0]; // @[LZD.scala 49:47]
  assign _T_191 = _T_184[0:0]; // @[LZD.scala 49:59]
  assign _T_192 = _T_185 ? _T_190 : _T_191; // @[LZD.scala 49:35]
  assign _T_194 = {_T_187,_T_189,_T_192}; // @[Cat.scala 29:58]
  assign _T_195 = _T_169[3:0]; // @[LZD.scala 44:32]
  assign _T_196 = _T_195[3:2]; // @[LZD.scala 43:32]
  assign _T_197 = _T_196 != 2'h0; // @[LZD.scala 39:14]
  assign _T_198 = _T_196[1]; // @[LZD.scala 39:21]
  assign _T_199 = _T_196[0]; // @[LZD.scala 39:30]
  assign _T_200 = ~ _T_199; // @[LZD.scala 39:27]
  assign _T_201 = _T_198 | _T_200; // @[LZD.scala 39:25]
  assign _T_202 = {_T_197,_T_201}; // @[Cat.scala 29:58]
  assign _T_203 = _T_195[1:0]; // @[LZD.scala 44:32]
  assign _T_204 = _T_203 != 2'h0; // @[LZD.scala 39:14]
  assign _T_205 = _T_203[1]; // @[LZD.scala 39:21]
  assign _T_206 = _T_203[0]; // @[LZD.scala 39:30]
  assign _T_207 = ~ _T_206; // @[LZD.scala 39:27]
  assign _T_208 = _T_205 | _T_207; // @[LZD.scala 39:25]
  assign _T_209 = {_T_204,_T_208}; // @[Cat.scala 29:58]
  assign _T_210 = _T_202[1]; // @[Shift.scala 12:21]
  assign _T_211 = _T_209[1]; // @[Shift.scala 12:21]
  assign _T_212 = _T_210 | _T_211; // @[LZD.scala 49:16]
  assign _T_213 = ~ _T_211; // @[LZD.scala 49:27]
  assign _T_214 = _T_210 | _T_213; // @[LZD.scala 49:25]
  assign _T_215 = _T_202[0:0]; // @[LZD.scala 49:47]
  assign _T_216 = _T_209[0:0]; // @[LZD.scala 49:59]
  assign _T_217 = _T_210 ? _T_215 : _T_216; // @[LZD.scala 49:35]
  assign _T_219 = {_T_212,_T_214,_T_217}; // @[Cat.scala 29:58]
  assign _T_220 = _T_194[2]; // @[Shift.scala 12:21]
  assign _T_221 = _T_219[2]; // @[Shift.scala 12:21]
  assign _T_222 = _T_220 | _T_221; // @[LZD.scala 49:16]
  assign _T_223 = ~ _T_221; // @[LZD.scala 49:27]
  assign _T_224 = _T_220 | _T_223; // @[LZD.scala 49:25]
  assign _T_225 = _T_194[1:0]; // @[LZD.scala 49:47]
  assign _T_226 = _T_219[1:0]; // @[LZD.scala 49:59]
  assign _T_227 = _T_220 ? _T_225 : _T_226; // @[LZD.scala 49:35]
  assign _T_229 = {_T_222,_T_224,_T_227}; // @[Cat.scala 29:58]
  assign _T_230 = _T_168[5:0]; // @[LZD.scala 44:32]
  assign _T_231 = _T_230[5:2]; // @[LZD.scala 43:32]
  assign _T_232 = _T_231[3:2]; // @[LZD.scala 43:32]
  assign _T_233 = _T_232 != 2'h0; // @[LZD.scala 39:14]
  assign _T_234 = _T_232[1]; // @[LZD.scala 39:21]
  assign _T_235 = _T_232[0]; // @[LZD.scala 39:30]
  assign _T_236 = ~ _T_235; // @[LZD.scala 39:27]
  assign _T_237 = _T_234 | _T_236; // @[LZD.scala 39:25]
  assign _T_238 = {_T_233,_T_237}; // @[Cat.scala 29:58]
  assign _T_239 = _T_231[1:0]; // @[LZD.scala 44:32]
  assign _T_240 = _T_239 != 2'h0; // @[LZD.scala 39:14]
  assign _T_241 = _T_239[1]; // @[LZD.scala 39:21]
  assign _T_242 = _T_239[0]; // @[LZD.scala 39:30]
  assign _T_243 = ~ _T_242; // @[LZD.scala 39:27]
  assign _T_244 = _T_241 | _T_243; // @[LZD.scala 39:25]
  assign _T_245 = {_T_240,_T_244}; // @[Cat.scala 29:58]
  assign _T_246 = _T_238[1]; // @[Shift.scala 12:21]
  assign _T_247 = _T_245[1]; // @[Shift.scala 12:21]
  assign _T_248 = _T_246 | _T_247; // @[LZD.scala 49:16]
  assign _T_249 = ~ _T_247; // @[LZD.scala 49:27]
  assign _T_250 = _T_246 | _T_249; // @[LZD.scala 49:25]
  assign _T_251 = _T_238[0:0]; // @[LZD.scala 49:47]
  assign _T_252 = _T_245[0:0]; // @[LZD.scala 49:59]
  assign _T_253 = _T_246 ? _T_251 : _T_252; // @[LZD.scala 49:35]
  assign _T_255 = {_T_248,_T_250,_T_253}; // @[Cat.scala 29:58]
  assign _T_256 = _T_230[1:0]; // @[LZD.scala 44:32]
  assign _T_257 = _T_256 != 2'h0; // @[LZD.scala 39:14]
  assign _T_258 = _T_256[1]; // @[LZD.scala 39:21]
  assign _T_259 = _T_256[0]; // @[LZD.scala 39:30]
  assign _T_260 = ~ _T_259; // @[LZD.scala 39:27]
  assign _T_261 = _T_258 | _T_260; // @[LZD.scala 39:25]
  assign _T_262 = {_T_257,_T_261}; // @[Cat.scala 29:58]
  assign _T_263 = _T_255[2]; // @[Shift.scala 12:21]
  assign _T_265 = _T_255[1:0]; // @[LZD.scala 55:32]
  assign _T_266 = _T_263 ? _T_265 : _T_262; // @[LZD.scala 55:20]
  assign _T_267 = {_T_263,_T_266}; // @[Cat.scala 29:58]
  assign _T_268 = _T_229[3]; // @[Shift.scala 12:21]
  assign _T_270 = _T_229[2:0]; // @[LZD.scala 55:32]
  assign _T_271 = _T_268 ? _T_270 : _T_267; // @[LZD.scala 55:20]
  assign _T_272 = {_T_268,_T_271}; // @[Cat.scala 29:58]
  assign _T_273 = ~ _T_272; // @[convert.scala 21:22]
  assign _T_274 = io_B[12:0]; // @[convert.scala 22:36]
  assign _T_275 = _T_273 < 4'hd; // @[Shift.scala 16:24]
  assign _T_277 = _T_273[3]; // @[Shift.scala 12:21]
  assign _T_278 = _T_274[4:0]; // @[Shift.scala 64:52]
  assign _T_280 = {_T_278,8'h0}; // @[Cat.scala 29:58]
  assign _T_281 = _T_277 ? _T_280 : _T_274; // @[Shift.scala 64:27]
  assign _T_282 = _T_273[2:0]; // @[Shift.scala 66:70]
  assign _T_283 = _T_282[2]; // @[Shift.scala 12:21]
  assign _T_284 = _T_281[8:0]; // @[Shift.scala 64:52]
  assign _T_286 = {_T_284,4'h0}; // @[Cat.scala 29:58]
  assign _T_287 = _T_283 ? _T_286 : _T_281; // @[Shift.scala 64:27]
  assign _T_288 = _T_282[1:0]; // @[Shift.scala 66:70]
  assign _T_289 = _T_288[1]; // @[Shift.scala 12:21]
  assign _T_290 = _T_287[10:0]; // @[Shift.scala 64:52]
  assign _T_292 = {_T_290,2'h0}; // @[Cat.scala 29:58]
  assign _T_293 = _T_289 ? _T_292 : _T_287; // @[Shift.scala 64:27]
  assign _T_294 = _T_288[0:0]; // @[Shift.scala 66:70]
  assign _T_296 = _T_293[11:0]; // @[Shift.scala 64:52]
  assign _T_297 = {_T_296,1'h0}; // @[Cat.scala 29:58]
  assign _T_298 = _T_294 ? _T_297 : _T_293; // @[Shift.scala 64:27]
  assign _T_299 = _T_275 ? _T_298 : 13'h0; // @[Shift.scala 16:10]
  assign _T_300 = _T_299[12:10]; // @[convert.scala 23:34]
  assign decB_fraction = _T_299[9:0]; // @[convert.scala 24:34]
  assign _T_302 = _T_165 == 1'h0; // @[convert.scala 25:26]
  assign _T_304 = _T_165 ? _T_273 : _T_272; // @[convert.scala 25:42]
  assign _T_307 = ~ _T_300; // @[convert.scala 26:67]
  assign _T_308 = _T_163 ? _T_307 : _T_300; // @[convert.scala 26:51]
  assign _T_309 = {_T_302,_T_304,_T_308}; // @[Cat.scala 29:58]
  assign _T_311 = io_B[14:0]; // @[convert.scala 29:56]
  assign _T_312 = _T_311 != 15'h0; // @[convert.scala 29:60]
  assign _T_313 = ~ _T_312; // @[convert.scala 29:41]
  assign decB_isNaR = _T_163 & _T_313; // @[convert.scala 29:39]
  assign _T_316 = _T_163 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_316 & _T_313; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_309); // @[convert.scala 32:24]
  assign aGTb = $signed(decA_scale) > $signed(decB_scale); // @[PositAdder.scala 24:32]
  assign greaterSign = aGTb ? _T_1 : _T_163; // @[PositAdder.scala 25:24]
  assign smallerSign = aGTb ? _T_163 : _T_1; // @[PositAdder.scala 26:24]
  assign greaterExp = aGTb ? $signed(decA_scale) : $signed(decB_scale); // @[PositAdder.scala 27:24]
  assign smallerExp = aGTb ? $signed(decB_scale) : $signed(decA_scale); // @[PositAdder.scala 28:24]
  assign greaterFrac = aGTb ? decA_fraction : decB_fraction; // @[PositAdder.scala 29:24]
  assign smallerFrac = aGTb ? decB_fraction : decA_fraction; // @[PositAdder.scala 30:24]
  assign smallerZero = aGTb ? decB_isZero : decA_isZero; // @[PositAdder.scala 31:24]
  assign _T_325 = $signed(greaterExp) - $signed(smallerExp); // @[PositAdder.scala 32:32]
  assign scale_diff = $signed(_T_325); // @[PositAdder.scala 32:32]
  assign _T_326 = ~ greaterSign; // @[PositAdder.scala 33:38]
  assign greaterSig = {greaterSign,_T_326,greaterFrac}; // @[Cat.scala 29:58]
  assign _T_328 = smallerSign | smallerZero; // @[PositAdder.scala 34:52]
  assign _T_329 = ~ _T_328; // @[PositAdder.scala 34:38]
  assign _T_332 = {smallerSign,_T_329,smallerFrac,3'h0}; // @[Cat.scala 29:58]
  assign _T_333 = $unsigned(scale_diff); // @[PositAdder.scala 35:68]
  assign _T_334 = _T_333 < 8'hf; // @[Shift.scala 39:24]
  assign _T_335 = _T_333[3:0]; // @[Shift.scala 40:44]
  assign _T_336 = _T_332[14:8]; // @[Shift.scala 90:30]
  assign _T_337 = _T_332[7:0]; // @[Shift.scala 90:48]
  assign _T_338 = _T_337 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_0 = {{6'd0}, _T_338}; // @[Shift.scala 90:39]
  assign _T_339 = _T_336 | _GEN_0; // @[Shift.scala 90:39]
  assign _T_340 = _T_335[3]; // @[Shift.scala 12:21]
  assign _T_341 = _T_332[14]; // @[Shift.scala 12:21]
  assign _T_343 = _T_341 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_344 = {_T_343,_T_339}; // @[Cat.scala 29:58]
  assign _T_345 = _T_340 ? _T_344 : _T_332; // @[Shift.scala 91:22]
  assign _T_346 = _T_335[2:0]; // @[Shift.scala 92:77]
  assign _T_347 = _T_345[14:4]; // @[Shift.scala 90:30]
  assign _T_348 = _T_345[3:0]; // @[Shift.scala 90:48]
  assign _T_349 = _T_348 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_1 = {{10'd0}, _T_349}; // @[Shift.scala 90:39]
  assign _T_350 = _T_347 | _GEN_1; // @[Shift.scala 90:39]
  assign _T_351 = _T_346[2]; // @[Shift.scala 12:21]
  assign _T_352 = _T_345[14]; // @[Shift.scala 12:21]
  assign _T_354 = _T_352 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_355 = {_T_354,_T_350}; // @[Cat.scala 29:58]
  assign _T_356 = _T_351 ? _T_355 : _T_345; // @[Shift.scala 91:22]
  assign _T_357 = _T_346[1:0]; // @[Shift.scala 92:77]
  assign _T_358 = _T_356[14:2]; // @[Shift.scala 90:30]
  assign _T_359 = _T_356[1:0]; // @[Shift.scala 90:48]
  assign _T_360 = _T_359 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_2 = {{12'd0}, _T_360}; // @[Shift.scala 90:39]
  assign _T_361 = _T_358 | _GEN_2; // @[Shift.scala 90:39]
  assign _T_362 = _T_357[1]; // @[Shift.scala 12:21]
  assign _T_363 = _T_356[14]; // @[Shift.scala 12:21]
  assign _T_365 = _T_363 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_366 = {_T_365,_T_361}; // @[Cat.scala 29:58]
  assign _T_367 = _T_362 ? _T_366 : _T_356; // @[Shift.scala 91:22]
  assign _T_368 = _T_357[0:0]; // @[Shift.scala 92:77]
  assign _T_369 = _T_367[14:1]; // @[Shift.scala 90:30]
  assign _T_370 = _T_367[0:0]; // @[Shift.scala 90:48]
  assign _GEN_3 = {{13'd0}, _T_370}; // @[Shift.scala 90:39]
  assign _T_372 = _T_369 | _GEN_3; // @[Shift.scala 90:39]
  assign _T_374 = _T_367[14]; // @[Shift.scala 12:21]
  assign _T_375 = {_T_374,_T_372}; // @[Cat.scala 29:58]
  assign _T_376 = _T_368 ? _T_375 : _T_367; // @[Shift.scala 91:22]
  assign _T_379 = _T_341 ? 15'h7fff : 15'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_334 ? _T_376 : _T_379; // @[Shift.scala 39:10]
  assign _T_380 = smallerSig[14:3]; // @[PositAdder.scala 36:45]
  assign rawSumSig = greaterSig + _T_380; // @[PositAdder.scala 36:32]
  assign _T_381 = _T_1 ^ _T_163; // @[PositAdder.scala 37:31]
  assign _T_382 = rawSumSig[12:12]; // @[PositAdder.scala 37:59]
  assign sumSign = _T_381 ^ _T_382; // @[PositAdder.scala 37:43]
  assign _T_383 = greaterSig + _T_380; // @[PositAdder.scala 38:48]
  assign _T_384 = smallerSig[2:0]; // @[PositAdder.scala 38:63]
  assign signSumSig = {sumSign,_T_383,_T_384}; // @[Cat.scala 29:58]
  assign _T_386 = signSumSig[15:1]; // @[PositAdder.scala 40:31]
  assign _T_387 = signSumSig[14:0]; // @[PositAdder.scala 40:66]
  assign sumXor = _T_386 ^ _T_387; // @[PositAdder.scala 40:49]
  assign _T_388 = sumXor[14:7]; // @[LZD.scala 43:32]
  assign _T_389 = _T_388[7:4]; // @[LZD.scala 43:32]
  assign _T_390 = _T_389[3:2]; // @[LZD.scala 43:32]
  assign _T_391 = _T_390 != 2'h0; // @[LZD.scala 39:14]
  assign _T_392 = _T_390[1]; // @[LZD.scala 39:21]
  assign _T_393 = _T_390[0]; // @[LZD.scala 39:30]
  assign _T_394 = ~ _T_393; // @[LZD.scala 39:27]
  assign _T_395 = _T_392 | _T_394; // @[LZD.scala 39:25]
  assign _T_396 = {_T_391,_T_395}; // @[Cat.scala 29:58]
  assign _T_397 = _T_389[1:0]; // @[LZD.scala 44:32]
  assign _T_398 = _T_397 != 2'h0; // @[LZD.scala 39:14]
  assign _T_399 = _T_397[1]; // @[LZD.scala 39:21]
  assign _T_400 = _T_397[0]; // @[LZD.scala 39:30]
  assign _T_401 = ~ _T_400; // @[LZD.scala 39:27]
  assign _T_402 = _T_399 | _T_401; // @[LZD.scala 39:25]
  assign _T_403 = {_T_398,_T_402}; // @[Cat.scala 29:58]
  assign _T_404 = _T_396[1]; // @[Shift.scala 12:21]
  assign _T_405 = _T_403[1]; // @[Shift.scala 12:21]
  assign _T_406 = _T_404 | _T_405; // @[LZD.scala 49:16]
  assign _T_407 = ~ _T_405; // @[LZD.scala 49:27]
  assign _T_408 = _T_404 | _T_407; // @[LZD.scala 49:25]
  assign _T_409 = _T_396[0:0]; // @[LZD.scala 49:47]
  assign _T_410 = _T_403[0:0]; // @[LZD.scala 49:59]
  assign _T_411 = _T_404 ? _T_409 : _T_410; // @[LZD.scala 49:35]
  assign _T_413 = {_T_406,_T_408,_T_411}; // @[Cat.scala 29:58]
  assign _T_414 = _T_388[3:0]; // @[LZD.scala 44:32]
  assign _T_415 = _T_414[3:2]; // @[LZD.scala 43:32]
  assign _T_416 = _T_415 != 2'h0; // @[LZD.scala 39:14]
  assign _T_417 = _T_415[1]; // @[LZD.scala 39:21]
  assign _T_418 = _T_415[0]; // @[LZD.scala 39:30]
  assign _T_419 = ~ _T_418; // @[LZD.scala 39:27]
  assign _T_420 = _T_417 | _T_419; // @[LZD.scala 39:25]
  assign _T_421 = {_T_416,_T_420}; // @[Cat.scala 29:58]
  assign _T_422 = _T_414[1:0]; // @[LZD.scala 44:32]
  assign _T_423 = _T_422 != 2'h0; // @[LZD.scala 39:14]
  assign _T_424 = _T_422[1]; // @[LZD.scala 39:21]
  assign _T_425 = _T_422[0]; // @[LZD.scala 39:30]
  assign _T_426 = ~ _T_425; // @[LZD.scala 39:27]
  assign _T_427 = _T_424 | _T_426; // @[LZD.scala 39:25]
  assign _T_428 = {_T_423,_T_427}; // @[Cat.scala 29:58]
  assign _T_429 = _T_421[1]; // @[Shift.scala 12:21]
  assign _T_430 = _T_428[1]; // @[Shift.scala 12:21]
  assign _T_431 = _T_429 | _T_430; // @[LZD.scala 49:16]
  assign _T_432 = ~ _T_430; // @[LZD.scala 49:27]
  assign _T_433 = _T_429 | _T_432; // @[LZD.scala 49:25]
  assign _T_434 = _T_421[0:0]; // @[LZD.scala 49:47]
  assign _T_435 = _T_428[0:0]; // @[LZD.scala 49:59]
  assign _T_436 = _T_429 ? _T_434 : _T_435; // @[LZD.scala 49:35]
  assign _T_438 = {_T_431,_T_433,_T_436}; // @[Cat.scala 29:58]
  assign _T_439 = _T_413[2]; // @[Shift.scala 12:21]
  assign _T_440 = _T_438[2]; // @[Shift.scala 12:21]
  assign _T_441 = _T_439 | _T_440; // @[LZD.scala 49:16]
  assign _T_442 = ~ _T_440; // @[LZD.scala 49:27]
  assign _T_443 = _T_439 | _T_442; // @[LZD.scala 49:25]
  assign _T_444 = _T_413[1:0]; // @[LZD.scala 49:47]
  assign _T_445 = _T_438[1:0]; // @[LZD.scala 49:59]
  assign _T_446 = _T_439 ? _T_444 : _T_445; // @[LZD.scala 49:35]
  assign _T_448 = {_T_441,_T_443,_T_446}; // @[Cat.scala 29:58]
  assign _T_449 = sumXor[6:0]; // @[LZD.scala 44:32]
  assign _T_450 = _T_449[6:3]; // @[LZD.scala 43:32]
  assign _T_451 = _T_450[3:2]; // @[LZD.scala 43:32]
  assign _T_452 = _T_451 != 2'h0; // @[LZD.scala 39:14]
  assign _T_453 = _T_451[1]; // @[LZD.scala 39:21]
  assign _T_454 = _T_451[0]; // @[LZD.scala 39:30]
  assign _T_455 = ~ _T_454; // @[LZD.scala 39:27]
  assign _T_456 = _T_453 | _T_455; // @[LZD.scala 39:25]
  assign _T_457 = {_T_452,_T_456}; // @[Cat.scala 29:58]
  assign _T_458 = _T_450[1:0]; // @[LZD.scala 44:32]
  assign _T_459 = _T_458 != 2'h0; // @[LZD.scala 39:14]
  assign _T_460 = _T_458[1]; // @[LZD.scala 39:21]
  assign _T_461 = _T_458[0]; // @[LZD.scala 39:30]
  assign _T_462 = ~ _T_461; // @[LZD.scala 39:27]
  assign _T_463 = _T_460 | _T_462; // @[LZD.scala 39:25]
  assign _T_464 = {_T_459,_T_463}; // @[Cat.scala 29:58]
  assign _T_465 = _T_457[1]; // @[Shift.scala 12:21]
  assign _T_466 = _T_464[1]; // @[Shift.scala 12:21]
  assign _T_467 = _T_465 | _T_466; // @[LZD.scala 49:16]
  assign _T_468 = ~ _T_466; // @[LZD.scala 49:27]
  assign _T_469 = _T_465 | _T_468; // @[LZD.scala 49:25]
  assign _T_470 = _T_457[0:0]; // @[LZD.scala 49:47]
  assign _T_471 = _T_464[0:0]; // @[LZD.scala 49:59]
  assign _T_472 = _T_465 ? _T_470 : _T_471; // @[LZD.scala 49:35]
  assign _T_474 = {_T_467,_T_469,_T_472}; // @[Cat.scala 29:58]
  assign _T_475 = _T_449[2:0]; // @[LZD.scala 44:32]
  assign _T_476 = _T_475[2:1]; // @[LZD.scala 43:32]
  assign _T_477 = _T_476 != 2'h0; // @[LZD.scala 39:14]
  assign _T_478 = _T_476[1]; // @[LZD.scala 39:21]
  assign _T_479 = _T_476[0]; // @[LZD.scala 39:30]
  assign _T_480 = ~ _T_479; // @[LZD.scala 39:27]
  assign _T_481 = _T_478 | _T_480; // @[LZD.scala 39:25]
  assign _T_482 = {_T_477,_T_481}; // @[Cat.scala 29:58]
  assign _T_483 = _T_475[0:0]; // @[LZD.scala 44:32]
  assign _T_485 = _T_482[1]; // @[Shift.scala 12:21]
  assign _T_487 = _T_482[0:0]; // @[LZD.scala 55:32]
  assign _T_488 = _T_485 ? _T_487 : _T_483; // @[LZD.scala 55:20]
  assign _T_489 = {_T_485,_T_488}; // @[Cat.scala 29:58]
  assign _T_490 = _T_474[2]; // @[Shift.scala 12:21]
  assign _T_492 = _T_474[1:0]; // @[LZD.scala 55:32]
  assign _T_493 = _T_490 ? _T_492 : _T_489; // @[LZD.scala 55:20]
  assign _T_494 = {_T_490,_T_493}; // @[Cat.scala 29:58]
  assign _T_495 = _T_448[3]; // @[Shift.scala 12:21]
  assign _T_497 = _T_448[2:0]; // @[LZD.scala 55:32]
  assign _T_498 = _T_495 ? _T_497 : _T_494; // @[LZD.scala 55:20]
  assign sumLZD = {_T_495,_T_498}; // @[Cat.scala 29:58]
  assign _T_499 = {1'h1,_T_495,_T_498}; // @[Cat.scala 29:58]
  assign _T_500 = $signed(_T_499); // @[PositAdder.scala 42:38]
  assign _T_502 = $signed(_T_500) + $signed(5'sh2); // @[PositAdder.scala 42:45]
  assign scaleBias = $signed(_T_502); // @[PositAdder.scala 42:45]
  assign _GEN_4 = {{3{scaleBias[4]}},scaleBias}; // @[PositAdder.scala 43:32]
  assign sumScale = $signed(greaterExp) + $signed(_GEN_4); // @[PositAdder.scala 43:32]
  assign overflow = $signed(sumScale) > $signed(9'sh70); // @[PositAdder.scala 44:30]
  assign normalShift = ~ sumLZD; // @[PositAdder.scala 45:22]
  assign _T_503 = signSumSig[13:0]; // @[PositAdder.scala 46:36]
  assign _T_504 = normalShift < 4'he; // @[Shift.scala 16:24]
  assign _T_506 = normalShift[3]; // @[Shift.scala 12:21]
  assign _T_507 = _T_503[5:0]; // @[Shift.scala 64:52]
  assign _T_509 = {_T_507,8'h0}; // @[Cat.scala 29:58]
  assign _T_510 = _T_506 ? _T_509 : _T_503; // @[Shift.scala 64:27]
  assign _T_511 = normalShift[2:0]; // @[Shift.scala 66:70]
  assign _T_512 = _T_511[2]; // @[Shift.scala 12:21]
  assign _T_513 = _T_510[9:0]; // @[Shift.scala 64:52]
  assign _T_515 = {_T_513,4'h0}; // @[Cat.scala 29:58]
  assign _T_516 = _T_512 ? _T_515 : _T_510; // @[Shift.scala 64:27]
  assign _T_517 = _T_511[1:0]; // @[Shift.scala 66:70]
  assign _T_518 = _T_517[1]; // @[Shift.scala 12:21]
  assign _T_519 = _T_516[11:0]; // @[Shift.scala 64:52]
  assign _T_521 = {_T_519,2'h0}; // @[Cat.scala 29:58]
  assign _T_522 = _T_518 ? _T_521 : _T_516; // @[Shift.scala 64:27]
  assign _T_523 = _T_517[0:0]; // @[Shift.scala 66:70]
  assign _T_525 = _T_522[12:0]; // @[Shift.scala 64:52]
  assign _T_526 = {_T_525,1'h0}; // @[Cat.scala 29:58]
  assign _T_527 = _T_523 ? _T_526 : _T_522; // @[Shift.scala 64:27]
  assign shiftSig = _T_504 ? _T_527 : 14'h0; // @[Shift.scala 16:10]
  assign _T_528 = overflow ? $signed(9'sh70) : $signed(sumScale); // @[PositAdder.scala 51:24]
  assign decS_fraction = shiftSig[13:4]; // @[PositAdder.scala 52:34]
  assign decS_isNaR = decA_isNaR | decB_isNaR; // @[PositAdder.scala 53:32]
  assign _T_531 = signSumSig != 16'h0; // @[PositAdder.scala 54:33]
  assign _T_532 = ~ _T_531; // @[PositAdder.scala 54:21]
  assign _T_533 = decA_isZero & decB_isZero; // @[PositAdder.scala 54:52]
  assign decS_isZero = _T_532 | _T_533; // @[PositAdder.scala 54:37]
  assign _T_535 = shiftSig[3:2]; // @[PositAdder.scala 55:33]
  assign _T_536 = shiftSig[1]; // @[PositAdder.scala 55:49]
  assign _T_537 = shiftSig[0]; // @[PositAdder.scala 55:63]
  assign _T_538 = _T_536 | _T_537; // @[PositAdder.scala 55:53]
  assign _GEN_5 = _T_528[7:0]; // @[PositAdder.scala 48:25 PositAdder.scala 51:18]
  assign decS_scale = $signed(_GEN_5); // @[PositAdder.scala 48:25 PositAdder.scala 51:18]
  assign _T_541 = decS_scale[2:0]; // @[convert.scala 46:61]
  assign _T_542 = ~ _T_541; // @[convert.scala 46:52]
  assign _T_544 = sumSign ? _T_542 : _T_541; // @[convert.scala 46:42]
  assign _T_545 = decS_scale[7:3]; // @[convert.scala 48:34]
  assign _T_546 = _T_545[4:4]; // @[convert.scala 49:36]
  assign _T_548 = ~ _T_545; // @[convert.scala 50:36]
  assign _T_549 = $signed(_T_548); // @[convert.scala 50:36]
  assign _T_550 = _T_546 ? $signed(_T_549) : $signed(_T_545); // @[convert.scala 50:28]
  assign _T_551 = _T_546 ^ sumSign; // @[convert.scala 51:31]
  assign _T_552 = ~ _T_551; // @[convert.scala 52:43]
  assign _T_556 = {_T_552,_T_551,_T_544,decS_fraction,_T_535,_T_538}; // @[Cat.scala 29:58]
  assign _T_557 = $unsigned(_T_550); // @[Shift.scala 39:17]
  assign _T_558 = _T_557 < 5'h12; // @[Shift.scala 39:24]
  assign _T_560 = _T_556[17:16]; // @[Shift.scala 90:30]
  assign _T_561 = _T_556[15:0]; // @[Shift.scala 90:48]
  assign _T_562 = _T_561 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_6 = {{1'd0}, _T_562}; // @[Shift.scala 90:39]
  assign _T_563 = _T_560 | _GEN_6; // @[Shift.scala 90:39]
  assign _T_564 = _T_557[4]; // @[Shift.scala 12:21]
  assign _T_565 = _T_556[17]; // @[Shift.scala 12:21]
  assign _T_567 = _T_565 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_568 = {_T_567,_T_563}; // @[Cat.scala 29:58]
  assign _T_569 = _T_564 ? _T_568 : _T_556; // @[Shift.scala 91:22]
  assign _T_570 = _T_557[3:0]; // @[Shift.scala 92:77]
  assign _T_571 = _T_569[17:8]; // @[Shift.scala 90:30]
  assign _T_572 = _T_569[7:0]; // @[Shift.scala 90:48]
  assign _T_573 = _T_572 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_7 = {{9'd0}, _T_573}; // @[Shift.scala 90:39]
  assign _T_574 = _T_571 | _GEN_7; // @[Shift.scala 90:39]
  assign _T_575 = _T_570[3]; // @[Shift.scala 12:21]
  assign _T_576 = _T_569[17]; // @[Shift.scala 12:21]
  assign _T_578 = _T_576 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_579 = {_T_578,_T_574}; // @[Cat.scala 29:58]
  assign _T_580 = _T_575 ? _T_579 : _T_569; // @[Shift.scala 91:22]
  assign _T_581 = _T_570[2:0]; // @[Shift.scala 92:77]
  assign _T_582 = _T_580[17:4]; // @[Shift.scala 90:30]
  assign _T_583 = _T_580[3:0]; // @[Shift.scala 90:48]
  assign _T_584 = _T_583 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_8 = {{13'd0}, _T_584}; // @[Shift.scala 90:39]
  assign _T_585 = _T_582 | _GEN_8; // @[Shift.scala 90:39]
  assign _T_586 = _T_581[2]; // @[Shift.scala 12:21]
  assign _T_587 = _T_580[17]; // @[Shift.scala 12:21]
  assign _T_589 = _T_587 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_590 = {_T_589,_T_585}; // @[Cat.scala 29:58]
  assign _T_591 = _T_586 ? _T_590 : _T_580; // @[Shift.scala 91:22]
  assign _T_592 = _T_581[1:0]; // @[Shift.scala 92:77]
  assign _T_593 = _T_591[17:2]; // @[Shift.scala 90:30]
  assign _T_594 = _T_591[1:0]; // @[Shift.scala 90:48]
  assign _T_595 = _T_594 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_9 = {{15'd0}, _T_595}; // @[Shift.scala 90:39]
  assign _T_596 = _T_593 | _GEN_9; // @[Shift.scala 90:39]
  assign _T_597 = _T_592[1]; // @[Shift.scala 12:21]
  assign _T_598 = _T_591[17]; // @[Shift.scala 12:21]
  assign _T_600 = _T_598 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_601 = {_T_600,_T_596}; // @[Cat.scala 29:58]
  assign _T_602 = _T_597 ? _T_601 : _T_591; // @[Shift.scala 91:22]
  assign _T_603 = _T_592[0:0]; // @[Shift.scala 92:77]
  assign _T_604 = _T_602[17:1]; // @[Shift.scala 90:30]
  assign _T_605 = _T_602[0:0]; // @[Shift.scala 90:48]
  assign _GEN_10 = {{16'd0}, _T_605}; // @[Shift.scala 90:39]
  assign _T_607 = _T_604 | _GEN_10; // @[Shift.scala 90:39]
  assign _T_609 = _T_602[17]; // @[Shift.scala 12:21]
  assign _T_610 = {_T_609,_T_607}; // @[Cat.scala 29:58]
  assign _T_611 = _T_603 ? _T_610 : _T_602; // @[Shift.scala 91:22]
  assign _T_614 = _T_565 ? 18'h3ffff : 18'h0; // @[Bitwise.scala 71:12]
  assign _T_615 = _T_558 ? _T_611 : _T_614; // @[Shift.scala 39:10]
  assign _T_616 = _T_615[3]; // @[convert.scala 55:31]
  assign _T_617 = _T_615[2]; // @[convert.scala 56:31]
  assign _T_618 = _T_615[1]; // @[convert.scala 57:31]
  assign _T_619 = _T_615[0]; // @[convert.scala 58:31]
  assign _T_620 = _T_615[17:3]; // @[convert.scala 59:69]
  assign _T_621 = _T_620 != 15'h0; // @[convert.scala 59:81]
  assign _T_622 = ~ _T_621; // @[convert.scala 59:50]
  assign _T_624 = _T_620 == 15'h7fff; // @[convert.scala 60:81]
  assign _T_625 = _T_616 | _T_618; // @[convert.scala 61:44]
  assign _T_626 = _T_625 | _T_619; // @[convert.scala 61:52]
  assign _T_627 = _T_617 & _T_626; // @[convert.scala 61:36]
  assign _T_628 = ~ _T_624; // @[convert.scala 62:63]
  assign _T_629 = _T_628 & _T_627; // @[convert.scala 62:103]
  assign _T_630 = _T_622 | _T_629; // @[convert.scala 62:60]
  assign _GEN_11 = {{14'd0}, _T_630}; // @[convert.scala 63:56]
  assign _T_633 = _T_620 + _GEN_11; // @[convert.scala 63:56]
  assign _T_634 = {sumSign,_T_633}; // @[Cat.scala 29:58]
  assign _T_636 = decS_isZero ? 16'h0 : _T_634; // @[Mux.scala 87:16]
  assign io_S = decS_isNaR ? 16'h8000 : _T_636; // @[PositAdder.scala 57:8]
endmodule
