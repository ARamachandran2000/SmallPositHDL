module PositFMA8_2(
  input        clock,
  input        reset,
  input        io_inValid,
  input  [1:0] io_fmaOp,
  input  [7:0] io_A,
  input  [7:0] io_B,
  input  [7:0] io_C,
  output [7:0] io_F,
  output       io_outValid
);
  wire  _T; // @[PositFMA.scala 47:36]
  wire [7:0] _T_2; // @[Bitwise.scala 71:12]
  wire [7:0] _T_3; // @[PositFMA.scala 47:41]
  wire [7:0] _GEN_10; // @[PositFMA.scala 47:49]
  wire [7:0] realA; // @[PositFMA.scala 47:49]
  wire  _T_6; // @[PositFMA.scala 48:36]
  wire [7:0] _T_8; // @[Bitwise.scala 71:12]
  wire [7:0] _T_9; // @[PositFMA.scala 48:41]
  wire [7:0] _GEN_11; // @[PositFMA.scala 48:49]
  wire [7:0] realC; // @[PositFMA.scala 48:49]
  wire  _T_13; // @[convert.scala 18:24]
  wire  _T_14; // @[convert.scala 18:40]
  wire  _T_15; // @[convert.scala 18:36]
  wire [5:0] _T_16; // @[convert.scala 19:24]
  wire [5:0] _T_17; // @[convert.scala 19:43]
  wire [5:0] _T_18; // @[convert.scala 19:39]
  wire [3:0] _T_19; // @[LZD.scala 43:32]
  wire [1:0] _T_20; // @[LZD.scala 43:32]
  wire  _T_21; // @[LZD.scala 39:14]
  wire  _T_22; // @[LZD.scala 39:21]
  wire  _T_23; // @[LZD.scala 39:30]
  wire  _T_24; // @[LZD.scala 39:27]
  wire  _T_25; // @[LZD.scala 39:25]
  wire [1:0] _T_26; // @[Cat.scala 29:58]
  wire [1:0] _T_27; // @[LZD.scala 44:32]
  wire  _T_28; // @[LZD.scala 39:14]
  wire  _T_29; // @[LZD.scala 39:21]
  wire  _T_30; // @[LZD.scala 39:30]
  wire  _T_31; // @[LZD.scala 39:27]
  wire  _T_32; // @[LZD.scala 39:25]
  wire [1:0] _T_33; // @[Cat.scala 29:58]
  wire  _T_34; // @[Shift.scala 12:21]
  wire  _T_35; // @[Shift.scala 12:21]
  wire  _T_36; // @[LZD.scala 49:16]
  wire  _T_37; // @[LZD.scala 49:27]
  wire  _T_38; // @[LZD.scala 49:25]
  wire  _T_39; // @[LZD.scala 49:47]
  wire  _T_40; // @[LZD.scala 49:59]
  wire  _T_41; // @[LZD.scala 49:35]
  wire [2:0] _T_43; // @[Cat.scala 29:58]
  wire [1:0] _T_44; // @[LZD.scala 44:32]
  wire  _T_45; // @[LZD.scala 39:14]
  wire  _T_46; // @[LZD.scala 39:21]
  wire  _T_47; // @[LZD.scala 39:30]
  wire  _T_48; // @[LZD.scala 39:27]
  wire  _T_49; // @[LZD.scala 39:25]
  wire [1:0] _T_50; // @[Cat.scala 29:58]
  wire  _T_51; // @[Shift.scala 12:21]
  wire [1:0] _T_53; // @[LZD.scala 55:32]
  wire [1:0] _T_54; // @[LZD.scala 55:20]
  wire [2:0] _T_55; // @[Cat.scala 29:58]
  wire [2:0] _T_56; // @[convert.scala 21:22]
  wire [4:0] _T_57; // @[convert.scala 22:36]
  wire  _T_58; // @[Shift.scala 16:24]
  wire  _T_60; // @[Shift.scala 12:21]
  wire  _T_61; // @[Shift.scala 64:52]
  wire [4:0] _T_63; // @[Cat.scala 29:58]
  wire [4:0] _T_64; // @[Shift.scala 64:27]
  wire [1:0] _T_65; // @[Shift.scala 66:70]
  wire  _T_66; // @[Shift.scala 12:21]
  wire [2:0] _T_67; // @[Shift.scala 64:52]
  wire [4:0] _T_69; // @[Cat.scala 29:58]
  wire [4:0] _T_70; // @[Shift.scala 64:27]
  wire  _T_71; // @[Shift.scala 66:70]
  wire [3:0] _T_73; // @[Shift.scala 64:52]
  wire [4:0] _T_74; // @[Cat.scala 29:58]
  wire [4:0] _T_75; // @[Shift.scala 64:27]
  wire [4:0] _T_76; // @[Shift.scala 16:10]
  wire [1:0] _T_77; // @[convert.scala 23:34]
  wire [2:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_79; // @[convert.scala 25:26]
  wire [2:0] _T_81; // @[convert.scala 25:42]
  wire [1:0] _T_84; // @[convert.scala 26:67]
  wire [1:0] _T_85; // @[convert.scala 26:51]
  wire [5:0] _T_86; // @[Cat.scala 29:58]
  wire [6:0] _T_88; // @[convert.scala 29:56]
  wire  _T_89; // @[convert.scala 29:60]
  wire  _T_90; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_93; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [5:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_102; // @[convert.scala 18:24]
  wire  _T_103; // @[convert.scala 18:40]
  wire  _T_104; // @[convert.scala 18:36]
  wire [5:0] _T_105; // @[convert.scala 19:24]
  wire [5:0] _T_106; // @[convert.scala 19:43]
  wire [5:0] _T_107; // @[convert.scala 19:39]
  wire [3:0] _T_108; // @[LZD.scala 43:32]
  wire [1:0] _T_109; // @[LZD.scala 43:32]
  wire  _T_110; // @[LZD.scala 39:14]
  wire  _T_111; // @[LZD.scala 39:21]
  wire  _T_112; // @[LZD.scala 39:30]
  wire  _T_113; // @[LZD.scala 39:27]
  wire  _T_114; // @[LZD.scala 39:25]
  wire [1:0] _T_115; // @[Cat.scala 29:58]
  wire [1:0] _T_116; // @[LZD.scala 44:32]
  wire  _T_117; // @[LZD.scala 39:14]
  wire  _T_118; // @[LZD.scala 39:21]
  wire  _T_119; // @[LZD.scala 39:30]
  wire  _T_120; // @[LZD.scala 39:27]
  wire  _T_121; // @[LZD.scala 39:25]
  wire [1:0] _T_122; // @[Cat.scala 29:58]
  wire  _T_123; // @[Shift.scala 12:21]
  wire  _T_124; // @[Shift.scala 12:21]
  wire  _T_125; // @[LZD.scala 49:16]
  wire  _T_126; // @[LZD.scala 49:27]
  wire  _T_127; // @[LZD.scala 49:25]
  wire  _T_128; // @[LZD.scala 49:47]
  wire  _T_129; // @[LZD.scala 49:59]
  wire  _T_130; // @[LZD.scala 49:35]
  wire [2:0] _T_132; // @[Cat.scala 29:58]
  wire [1:0] _T_133; // @[LZD.scala 44:32]
  wire  _T_134; // @[LZD.scala 39:14]
  wire  _T_135; // @[LZD.scala 39:21]
  wire  _T_136; // @[LZD.scala 39:30]
  wire  _T_137; // @[LZD.scala 39:27]
  wire  _T_138; // @[LZD.scala 39:25]
  wire [1:0] _T_139; // @[Cat.scala 29:58]
  wire  _T_140; // @[Shift.scala 12:21]
  wire [1:0] _T_142; // @[LZD.scala 55:32]
  wire [1:0] _T_143; // @[LZD.scala 55:20]
  wire [2:0] _T_144; // @[Cat.scala 29:58]
  wire [2:0] _T_145; // @[convert.scala 21:22]
  wire [4:0] _T_146; // @[convert.scala 22:36]
  wire  _T_147; // @[Shift.scala 16:24]
  wire  _T_149; // @[Shift.scala 12:21]
  wire  _T_150; // @[Shift.scala 64:52]
  wire [4:0] _T_152; // @[Cat.scala 29:58]
  wire [4:0] _T_153; // @[Shift.scala 64:27]
  wire [1:0] _T_154; // @[Shift.scala 66:70]
  wire  _T_155; // @[Shift.scala 12:21]
  wire [2:0] _T_156; // @[Shift.scala 64:52]
  wire [4:0] _T_158; // @[Cat.scala 29:58]
  wire [4:0] _T_159; // @[Shift.scala 64:27]
  wire  _T_160; // @[Shift.scala 66:70]
  wire [3:0] _T_162; // @[Shift.scala 64:52]
  wire [4:0] _T_163; // @[Cat.scala 29:58]
  wire [4:0] _T_164; // @[Shift.scala 64:27]
  wire [4:0] _T_165; // @[Shift.scala 16:10]
  wire [1:0] _T_166; // @[convert.scala 23:34]
  wire [2:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_168; // @[convert.scala 25:26]
  wire [2:0] _T_170; // @[convert.scala 25:42]
  wire [1:0] _T_173; // @[convert.scala 26:67]
  wire [1:0] _T_174; // @[convert.scala 26:51]
  wire [5:0] _T_175; // @[Cat.scala 29:58]
  wire [6:0] _T_177; // @[convert.scala 29:56]
  wire  _T_178; // @[convert.scala 29:60]
  wire  _T_179; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_182; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [5:0] decB_scale; // @[convert.scala 32:24]
  wire  _T_191; // @[convert.scala 18:24]
  wire  _T_192; // @[convert.scala 18:40]
  wire  _T_193; // @[convert.scala 18:36]
  wire [5:0] _T_194; // @[convert.scala 19:24]
  wire [5:0] _T_195; // @[convert.scala 19:43]
  wire [5:0] _T_196; // @[convert.scala 19:39]
  wire [3:0] _T_197; // @[LZD.scala 43:32]
  wire [1:0] _T_198; // @[LZD.scala 43:32]
  wire  _T_199; // @[LZD.scala 39:14]
  wire  _T_200; // @[LZD.scala 39:21]
  wire  _T_201; // @[LZD.scala 39:30]
  wire  _T_202; // @[LZD.scala 39:27]
  wire  _T_203; // @[LZD.scala 39:25]
  wire [1:0] _T_204; // @[Cat.scala 29:58]
  wire [1:0] _T_205; // @[LZD.scala 44:32]
  wire  _T_206; // @[LZD.scala 39:14]
  wire  _T_207; // @[LZD.scala 39:21]
  wire  _T_208; // @[LZD.scala 39:30]
  wire  _T_209; // @[LZD.scala 39:27]
  wire  _T_210; // @[LZD.scala 39:25]
  wire [1:0] _T_211; // @[Cat.scala 29:58]
  wire  _T_212; // @[Shift.scala 12:21]
  wire  _T_213; // @[Shift.scala 12:21]
  wire  _T_214; // @[LZD.scala 49:16]
  wire  _T_215; // @[LZD.scala 49:27]
  wire  _T_216; // @[LZD.scala 49:25]
  wire  _T_217; // @[LZD.scala 49:47]
  wire  _T_218; // @[LZD.scala 49:59]
  wire  _T_219; // @[LZD.scala 49:35]
  wire [2:0] _T_221; // @[Cat.scala 29:58]
  wire [1:0] _T_222; // @[LZD.scala 44:32]
  wire  _T_223; // @[LZD.scala 39:14]
  wire  _T_224; // @[LZD.scala 39:21]
  wire  _T_225; // @[LZD.scala 39:30]
  wire  _T_226; // @[LZD.scala 39:27]
  wire  _T_227; // @[LZD.scala 39:25]
  wire [1:0] _T_228; // @[Cat.scala 29:58]
  wire  _T_229; // @[Shift.scala 12:21]
  wire [1:0] _T_231; // @[LZD.scala 55:32]
  wire [1:0] _T_232; // @[LZD.scala 55:20]
  wire [2:0] _T_233; // @[Cat.scala 29:58]
  wire [2:0] _T_234; // @[convert.scala 21:22]
  wire [4:0] _T_235; // @[convert.scala 22:36]
  wire  _T_236; // @[Shift.scala 16:24]
  wire  _T_238; // @[Shift.scala 12:21]
  wire  _T_239; // @[Shift.scala 64:52]
  wire [4:0] _T_241; // @[Cat.scala 29:58]
  wire [4:0] _T_242; // @[Shift.scala 64:27]
  wire [1:0] _T_243; // @[Shift.scala 66:70]
  wire  _T_244; // @[Shift.scala 12:21]
  wire [2:0] _T_245; // @[Shift.scala 64:52]
  wire [4:0] _T_247; // @[Cat.scala 29:58]
  wire [4:0] _T_248; // @[Shift.scala 64:27]
  wire  _T_249; // @[Shift.scala 66:70]
  wire [3:0] _T_251; // @[Shift.scala 64:52]
  wire [4:0] _T_252; // @[Cat.scala 29:58]
  wire [4:0] _T_253; // @[Shift.scala 64:27]
  wire [4:0] _T_254; // @[Shift.scala 16:10]
  wire [1:0] _T_255; // @[convert.scala 23:34]
  wire [2:0] decC_fraction; // @[convert.scala 24:34]
  wire  _T_257; // @[convert.scala 25:26]
  wire [2:0] _T_259; // @[convert.scala 25:42]
  wire [1:0] _T_262; // @[convert.scala 26:67]
  wire [1:0] _T_263; // @[convert.scala 26:51]
  wire [5:0] _T_264; // @[Cat.scala 29:58]
  wire [6:0] _T_266; // @[convert.scala 29:56]
  wire  _T_267; // @[convert.scala 29:60]
  wire  _T_268; // @[convert.scala 29:41]
  wire  decC_isNaR; // @[convert.scala 29:39]
  wire  _T_271; // @[convert.scala 30:19]
  wire  decC_isZero; // @[convert.scala 30:41]
  wire [5:0] decC_scale; // @[convert.scala 32:24]
  wire  _T_279; // @[PositFMA.scala 58:30]
  wire  outIsNaR; // @[PositFMA.scala 58:44]
  wire  _T_280; // @[PositFMA.scala 59:34]
  wire  _T_281; // @[PositFMA.scala 59:47]
  wire  _T_282; // @[PositFMA.scala 59:45]
  wire [4:0] _T_284; // @[Cat.scala 29:58]
  wire [4:0] sigA; // @[PositFMA.scala 59:76]
  wire  _T_285; // @[PositFMA.scala 60:34]
  wire  _T_286; // @[PositFMA.scala 60:47]
  wire  _T_287; // @[PositFMA.scala 60:45]
  wire [4:0] _T_289; // @[Cat.scala 29:58]
  wire [4:0] sigB; // @[PositFMA.scala 60:76]
  wire [9:0] _T_290; // @[PositFMA.scala 61:25]
  wire [9:0] sigP; // @[PositFMA.scala 61:33]
  wire [1:0] head2; // @[PositFMA.scala 62:28]
  wire  _T_291; // @[PositFMA.scala 63:31]
  wire  _T_292; // @[PositFMA.scala 63:25]
  wire  _T_293; // @[PositFMA.scala 63:42]
  wire  addTwo; // @[PositFMA.scala 63:35]
  wire  _T_294; // @[PositFMA.scala 65:23]
  wire  _T_295; // @[PositFMA.scala 65:49]
  wire  addOne; // @[PositFMA.scala 65:43]
  wire [1:0] _T_296; // @[Cat.scala 29:58]
  wire [2:0] expBias; // @[PositFMA.scala 66:39]
  wire  mulSign; // @[PositFMA.scala 67:28]
  wire [6:0] _T_297; // @[PositFMA.scala 69:30]
  wire [6:0] _GEN_12; // @[PositFMA.scala 69:44]
  wire [6:0] _T_299; // @[PositFMA.scala 69:44]
  wire [6:0] mulScale; // @[PositFMA.scala 69:44]
  wire [7:0] _T_300; // @[PositFMA.scala 72:29]
  wire [6:0] _T_301; // @[PositFMA.scala 73:29]
  wire [7:0] _T_302; // @[PositFMA.scala 73:48]
  wire [7:0] mulSigTmp; // @[PositFMA.scala 70:22]
  wire  _T_304; // @[PositFMA.scala 77:39]
  wire  _T_305; // @[PositFMA.scala 77:43]
  wire [6:0] _T_306; // @[PositFMA.scala 78:39]
  wire [8:0] mulSig; // @[Cat.scala 29:58]
  reg  outIsNaR_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg [8:0] mulSig_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg [2:0] addFrac_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [6:0] mulScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [5:0] addScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  addSign_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  addZero_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  inValid_phase2; // @[Valid.scala 117:22]
  reg [31:0] _RAND_7;
  wire  _T_332; // @[PositFMA.scala 107:29]
  wire  _T_333; // @[PositFMA.scala 107:47]
  wire  _T_334; // @[PositFMA.scala 107:45]
  wire [8:0] extAddSig; // @[Cat.scala 29:58]
  wire [6:0] _GEN_13; // @[PositFMA.scala 111:39]
  wire  mulGreater; // @[PositFMA.scala 111:39]
  wire [6:0] greaterScale; // @[PositFMA.scala 112:26]
  wire [6:0] smallerScale; // @[PositFMA.scala 113:26]
  wire [6:0] _T_338; // @[PositFMA.scala 114:36]
  wire [6:0] scaleDiff; // @[PositFMA.scala 114:36]
  wire [8:0] greaterSig; // @[PositFMA.scala 115:26]
  wire [8:0] smallerSigTmp; // @[PositFMA.scala 116:26]
  wire [6:0] _T_339; // @[PositFMA.scala 117:69]
  wire  _T_340; // @[Shift.scala 39:24]
  wire [3:0] _T_341; // @[Shift.scala 40:44]
  wire  _T_342; // @[Shift.scala 90:30]
  wire [7:0] _T_343; // @[Shift.scala 90:48]
  wire  _T_344; // @[Shift.scala 90:57]
  wire  _T_345; // @[Shift.scala 90:39]
  wire  _T_346; // @[Shift.scala 12:21]
  wire  _T_347; // @[Shift.scala 12:21]
  wire [7:0] _T_349; // @[Bitwise.scala 71:12]
  wire [8:0] _T_350; // @[Cat.scala 29:58]
  wire [8:0] _T_351; // @[Shift.scala 91:22]
  wire [2:0] _T_352; // @[Shift.scala 92:77]
  wire [4:0] _T_353; // @[Shift.scala 90:30]
  wire [3:0] _T_354; // @[Shift.scala 90:48]
  wire  _T_355; // @[Shift.scala 90:57]
  wire [4:0] _GEN_14; // @[Shift.scala 90:39]
  wire [4:0] _T_356; // @[Shift.scala 90:39]
  wire  _T_357; // @[Shift.scala 12:21]
  wire  _T_358; // @[Shift.scala 12:21]
  wire [3:0] _T_360; // @[Bitwise.scala 71:12]
  wire [8:0] _T_361; // @[Cat.scala 29:58]
  wire [8:0] _T_362; // @[Shift.scala 91:22]
  wire [1:0] _T_363; // @[Shift.scala 92:77]
  wire [6:0] _T_364; // @[Shift.scala 90:30]
  wire [1:0] _T_365; // @[Shift.scala 90:48]
  wire  _T_366; // @[Shift.scala 90:57]
  wire [6:0] _GEN_15; // @[Shift.scala 90:39]
  wire [6:0] _T_367; // @[Shift.scala 90:39]
  wire  _T_368; // @[Shift.scala 12:21]
  wire  _T_369; // @[Shift.scala 12:21]
  wire [1:0] _T_371; // @[Bitwise.scala 71:12]
  wire [8:0] _T_372; // @[Cat.scala 29:58]
  wire [8:0] _T_373; // @[Shift.scala 91:22]
  wire  _T_374; // @[Shift.scala 92:77]
  wire [7:0] _T_375; // @[Shift.scala 90:30]
  wire  _T_376; // @[Shift.scala 90:48]
  wire [7:0] _GEN_16; // @[Shift.scala 90:39]
  wire [7:0] _T_378; // @[Shift.scala 90:39]
  wire  _T_380; // @[Shift.scala 12:21]
  wire [8:0] _T_381; // @[Cat.scala 29:58]
  wire [8:0] _T_382; // @[Shift.scala 91:22]
  wire [8:0] _T_385; // @[Bitwise.scala 71:12]
  wire [8:0] smallerSig; // @[Shift.scala 39:10]
  wire [9:0] rawSumSig; // @[PositFMA.scala 118:34]
  wire  _T_386; // @[PositFMA.scala 119:42]
  wire  _T_387; // @[PositFMA.scala 119:46]
  wire  _T_388; // @[PositFMA.scala 119:79]
  wire  sumSign; // @[PositFMA.scala 119:63]
  wire [8:0] _T_390; // @[PositFMA.scala 120:50]
  wire [9:0] signSumSig; // @[Cat.scala 29:58]
  wire [8:0] _T_391; // @[PositFMA.scala 124:33]
  wire [8:0] _T_392; // @[PositFMA.scala 124:68]
  wire [8:0] sumXor; // @[PositFMA.scala 124:51]
  wire [7:0] _T_393; // @[LZD.scala 43:32]
  wire [3:0] _T_394; // @[LZD.scala 43:32]
  wire [1:0] _T_395; // @[LZD.scala 43:32]
  wire  _T_396; // @[LZD.scala 39:14]
  wire  _T_397; // @[LZD.scala 39:21]
  wire  _T_398; // @[LZD.scala 39:30]
  wire  _T_399; // @[LZD.scala 39:27]
  wire  _T_400; // @[LZD.scala 39:25]
  wire [1:0] _T_401; // @[Cat.scala 29:58]
  wire [1:0] _T_402; // @[LZD.scala 44:32]
  wire  _T_403; // @[LZD.scala 39:14]
  wire  _T_404; // @[LZD.scala 39:21]
  wire  _T_405; // @[LZD.scala 39:30]
  wire  _T_406; // @[LZD.scala 39:27]
  wire  _T_407; // @[LZD.scala 39:25]
  wire [1:0] _T_408; // @[Cat.scala 29:58]
  wire  _T_409; // @[Shift.scala 12:21]
  wire  _T_410; // @[Shift.scala 12:21]
  wire  _T_411; // @[LZD.scala 49:16]
  wire  _T_412; // @[LZD.scala 49:27]
  wire  _T_413; // @[LZD.scala 49:25]
  wire  _T_414; // @[LZD.scala 49:47]
  wire  _T_415; // @[LZD.scala 49:59]
  wire  _T_416; // @[LZD.scala 49:35]
  wire [2:0] _T_418; // @[Cat.scala 29:58]
  wire [3:0] _T_419; // @[LZD.scala 44:32]
  wire [1:0] _T_420; // @[LZD.scala 43:32]
  wire  _T_421; // @[LZD.scala 39:14]
  wire  _T_422; // @[LZD.scala 39:21]
  wire  _T_423; // @[LZD.scala 39:30]
  wire  _T_424; // @[LZD.scala 39:27]
  wire  _T_425; // @[LZD.scala 39:25]
  wire [1:0] _T_426; // @[Cat.scala 29:58]
  wire [1:0] _T_427; // @[LZD.scala 44:32]
  wire  _T_428; // @[LZD.scala 39:14]
  wire  _T_429; // @[LZD.scala 39:21]
  wire  _T_430; // @[LZD.scala 39:30]
  wire  _T_431; // @[LZD.scala 39:27]
  wire  _T_432; // @[LZD.scala 39:25]
  wire [1:0] _T_433; // @[Cat.scala 29:58]
  wire  _T_434; // @[Shift.scala 12:21]
  wire  _T_435; // @[Shift.scala 12:21]
  wire  _T_436; // @[LZD.scala 49:16]
  wire  _T_437; // @[LZD.scala 49:27]
  wire  _T_438; // @[LZD.scala 49:25]
  wire  _T_439; // @[LZD.scala 49:47]
  wire  _T_440; // @[LZD.scala 49:59]
  wire  _T_441; // @[LZD.scala 49:35]
  wire [2:0] _T_443; // @[Cat.scala 29:58]
  wire  _T_444; // @[Shift.scala 12:21]
  wire  _T_445; // @[Shift.scala 12:21]
  wire  _T_446; // @[LZD.scala 49:16]
  wire  _T_447; // @[LZD.scala 49:27]
  wire  _T_448; // @[LZD.scala 49:25]
  wire [1:0] _T_449; // @[LZD.scala 49:47]
  wire [1:0] _T_450; // @[LZD.scala 49:59]
  wire [1:0] _T_451; // @[LZD.scala 49:35]
  wire [3:0] _T_453; // @[Cat.scala 29:58]
  wire  _T_454; // @[LZD.scala 44:32]
  wire  _T_456; // @[Shift.scala 12:21]
  wire [2:0] _T_459; // @[Cat.scala 29:58]
  wire [2:0] _T_460; // @[LZD.scala 55:32]
  wire [2:0] _T_461; // @[LZD.scala 55:20]
  wire [3:0] sumLZD; // @[Cat.scala 29:58]
  wire [3:0] shiftValue; // @[PositFMA.scala 126:24]
  wire [7:0] _T_462; // @[PositFMA.scala 127:38]
  wire  _T_463; // @[Shift.scala 16:24]
  wire [2:0] _T_464; // @[Shift.scala 17:37]
  wire  _T_465; // @[Shift.scala 12:21]
  wire [3:0] _T_466; // @[Shift.scala 64:52]
  wire [7:0] _T_468; // @[Cat.scala 29:58]
  wire [7:0] _T_469; // @[Shift.scala 64:27]
  wire [1:0] _T_470; // @[Shift.scala 66:70]
  wire  _T_471; // @[Shift.scala 12:21]
  wire [5:0] _T_472; // @[Shift.scala 64:52]
  wire [7:0] _T_474; // @[Cat.scala 29:58]
  wire [7:0] _T_475; // @[Shift.scala 64:27]
  wire  _T_476; // @[Shift.scala 66:70]
  wire [6:0] _T_478; // @[Shift.scala 64:52]
  wire [7:0] _T_479; // @[Cat.scala 29:58]
  wire [7:0] _T_480; // @[Shift.scala 64:27]
  wire [7:0] normalFracTmp; // @[Shift.scala 16:10]
  wire [6:0] _T_482; // @[PositFMA.scala 130:36]
  wire [6:0] _T_483; // @[PositFMA.scala 130:36]
  wire [4:0] _T_484; // @[Cat.scala 29:58]
  wire [4:0] _T_485; // @[PositFMA.scala 130:61]
  wire [6:0] _GEN_17; // @[PositFMA.scala 130:42]
  wire [6:0] _T_487; // @[PositFMA.scala 130:42]
  wire [6:0] sumScale; // @[PositFMA.scala 130:42]
  wire [2:0] sumFrac; // @[PositFMA.scala 131:41]
  wire [4:0] grsTmp; // @[PositFMA.scala 134:41]
  wire [1:0] _T_488; // @[PositFMA.scala 137:40]
  wire [2:0] _T_489; // @[PositFMA.scala 137:56]
  wire  _T_490; // @[PositFMA.scala 137:60]
  wire  underflow; // @[PositFMA.scala 144:32]
  wire  overflow; // @[PositFMA.scala 145:32]
  wire  _T_491; // @[PositFMA.scala 154:32]
  wire  decF_isZero; // @[PositFMA.scala 154:20]
  wire [6:0] _T_493; // @[Mux.scala 87:16]
  wire [6:0] _T_494; // @[Mux.scala 87:16]
  wire [5:0] _GEN_18; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  wire [5:0] decF_scale; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  wire [1:0] _T_495; // @[convert.scala 46:61]
  wire [1:0] _T_496; // @[convert.scala 46:52]
  wire [1:0] _T_498; // @[convert.scala 46:42]
  wire [3:0] _T_499; // @[convert.scala 48:34]
  wire  _T_500; // @[convert.scala 49:36]
  wire [3:0] _T_502; // @[convert.scala 50:36]
  wire [3:0] _T_503; // @[convert.scala 50:36]
  wire [3:0] _T_504; // @[convert.scala 50:28]
  wire  _T_505; // @[convert.scala 51:31]
  wire  _T_506; // @[convert.scala 52:43]
  wire [9:0] _T_510; // @[Cat.scala 29:58]
  wire [3:0] _T_511; // @[Shift.scala 39:17]
  wire  _T_512; // @[Shift.scala 39:24]
  wire [1:0] _T_514; // @[Shift.scala 90:30]
  wire [7:0] _T_515; // @[Shift.scala 90:48]
  wire  _T_516; // @[Shift.scala 90:57]
  wire [1:0] _GEN_19; // @[Shift.scala 90:39]
  wire [1:0] _T_517; // @[Shift.scala 90:39]
  wire  _T_518; // @[Shift.scala 12:21]
  wire  _T_519; // @[Shift.scala 12:21]
  wire [7:0] _T_521; // @[Bitwise.scala 71:12]
  wire [9:0] _T_522; // @[Cat.scala 29:58]
  wire [9:0] _T_523; // @[Shift.scala 91:22]
  wire [2:0] _T_524; // @[Shift.scala 92:77]
  wire [5:0] _T_525; // @[Shift.scala 90:30]
  wire [3:0] _T_526; // @[Shift.scala 90:48]
  wire  _T_527; // @[Shift.scala 90:57]
  wire [5:0] _GEN_20; // @[Shift.scala 90:39]
  wire [5:0] _T_528; // @[Shift.scala 90:39]
  wire  _T_529; // @[Shift.scala 12:21]
  wire  _T_530; // @[Shift.scala 12:21]
  wire [3:0] _T_532; // @[Bitwise.scala 71:12]
  wire [9:0] _T_533; // @[Cat.scala 29:58]
  wire [9:0] _T_534; // @[Shift.scala 91:22]
  wire [1:0] _T_535; // @[Shift.scala 92:77]
  wire [7:0] _T_536; // @[Shift.scala 90:30]
  wire [1:0] _T_537; // @[Shift.scala 90:48]
  wire  _T_538; // @[Shift.scala 90:57]
  wire [7:0] _GEN_21; // @[Shift.scala 90:39]
  wire [7:0] _T_539; // @[Shift.scala 90:39]
  wire  _T_540; // @[Shift.scala 12:21]
  wire  _T_541; // @[Shift.scala 12:21]
  wire [1:0] _T_543; // @[Bitwise.scala 71:12]
  wire [9:0] _T_544; // @[Cat.scala 29:58]
  wire [9:0] _T_545; // @[Shift.scala 91:22]
  wire  _T_546; // @[Shift.scala 92:77]
  wire [8:0] _T_547; // @[Shift.scala 90:30]
  wire  _T_548; // @[Shift.scala 90:48]
  wire [8:0] _GEN_22; // @[Shift.scala 90:39]
  wire [8:0] _T_550; // @[Shift.scala 90:39]
  wire  _T_552; // @[Shift.scala 12:21]
  wire [9:0] _T_553; // @[Cat.scala 29:58]
  wire [9:0] _T_554; // @[Shift.scala 91:22]
  wire [9:0] _T_557; // @[Bitwise.scala 71:12]
  wire [9:0] _T_558; // @[Shift.scala 39:10]
  wire  _T_559; // @[convert.scala 55:31]
  wire  _T_560; // @[convert.scala 56:31]
  wire  _T_561; // @[convert.scala 57:31]
  wire  _T_562; // @[convert.scala 58:31]
  wire [6:0] _T_563; // @[convert.scala 59:69]
  wire  _T_564; // @[convert.scala 59:81]
  wire  _T_565; // @[convert.scala 59:50]
  wire  _T_567; // @[convert.scala 60:81]
  wire  _T_568; // @[convert.scala 61:44]
  wire  _T_569; // @[convert.scala 61:52]
  wire  _T_570; // @[convert.scala 61:36]
  wire  _T_571; // @[convert.scala 62:63]
  wire  _T_572; // @[convert.scala 62:103]
  wire  _T_573; // @[convert.scala 62:60]
  wire [6:0] _GEN_23; // @[convert.scala 63:56]
  wire [6:0] _T_576; // @[convert.scala 63:56]
  wire [7:0] _T_577; // @[Cat.scala 29:58]
  reg  _T_581; // @[Valid.scala 117:22]
  reg [31:0] _RAND_8;
  reg [7:0] _T_585; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  assign _T = io_fmaOp[1]; // @[PositFMA.scala 47:36]
  assign _T_2 = _T ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_3 = _T_2 ^ io_A; // @[PositFMA.scala 47:41]
  assign _GEN_10 = {{7'd0}, _T}; // @[PositFMA.scala 47:49]
  assign realA = _T_3 + _GEN_10; // @[PositFMA.scala 47:49]
  assign _T_6 = io_fmaOp[0]; // @[PositFMA.scala 48:36]
  assign _T_8 = _T_6 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_9 = _T_8 ^ io_C; // @[PositFMA.scala 48:41]
  assign _GEN_11 = {{7'd0}, _T_6}; // @[PositFMA.scala 48:49]
  assign realC = _T_9 + _GEN_11; // @[PositFMA.scala 48:49]
  assign _T_13 = realA[7]; // @[convert.scala 18:24]
  assign _T_14 = realA[6]; // @[convert.scala 18:40]
  assign _T_15 = _T_13 ^ _T_14; // @[convert.scala 18:36]
  assign _T_16 = realA[6:1]; // @[convert.scala 19:24]
  assign _T_17 = realA[5:0]; // @[convert.scala 19:43]
  assign _T_18 = _T_16 ^ _T_17; // @[convert.scala 19:39]
  assign _T_19 = _T_18[5:2]; // @[LZD.scala 43:32]
  assign _T_20 = _T_19[3:2]; // @[LZD.scala 43:32]
  assign _T_21 = _T_20 != 2'h0; // @[LZD.scala 39:14]
  assign _T_22 = _T_20[1]; // @[LZD.scala 39:21]
  assign _T_23 = _T_20[0]; // @[LZD.scala 39:30]
  assign _T_24 = ~ _T_23; // @[LZD.scala 39:27]
  assign _T_25 = _T_22 | _T_24; // @[LZD.scala 39:25]
  assign _T_26 = {_T_21,_T_25}; // @[Cat.scala 29:58]
  assign _T_27 = _T_19[1:0]; // @[LZD.scala 44:32]
  assign _T_28 = _T_27 != 2'h0; // @[LZD.scala 39:14]
  assign _T_29 = _T_27[1]; // @[LZD.scala 39:21]
  assign _T_30 = _T_27[0]; // @[LZD.scala 39:30]
  assign _T_31 = ~ _T_30; // @[LZD.scala 39:27]
  assign _T_32 = _T_29 | _T_31; // @[LZD.scala 39:25]
  assign _T_33 = {_T_28,_T_32}; // @[Cat.scala 29:58]
  assign _T_34 = _T_26[1]; // @[Shift.scala 12:21]
  assign _T_35 = _T_33[1]; // @[Shift.scala 12:21]
  assign _T_36 = _T_34 | _T_35; // @[LZD.scala 49:16]
  assign _T_37 = ~ _T_35; // @[LZD.scala 49:27]
  assign _T_38 = _T_34 | _T_37; // @[LZD.scala 49:25]
  assign _T_39 = _T_26[0:0]; // @[LZD.scala 49:47]
  assign _T_40 = _T_33[0:0]; // @[LZD.scala 49:59]
  assign _T_41 = _T_34 ? _T_39 : _T_40; // @[LZD.scala 49:35]
  assign _T_43 = {_T_36,_T_38,_T_41}; // @[Cat.scala 29:58]
  assign _T_44 = _T_18[1:0]; // @[LZD.scala 44:32]
  assign _T_45 = _T_44 != 2'h0; // @[LZD.scala 39:14]
  assign _T_46 = _T_44[1]; // @[LZD.scala 39:21]
  assign _T_47 = _T_44[0]; // @[LZD.scala 39:30]
  assign _T_48 = ~ _T_47; // @[LZD.scala 39:27]
  assign _T_49 = _T_46 | _T_48; // @[LZD.scala 39:25]
  assign _T_50 = {_T_45,_T_49}; // @[Cat.scala 29:58]
  assign _T_51 = _T_43[2]; // @[Shift.scala 12:21]
  assign _T_53 = _T_43[1:0]; // @[LZD.scala 55:32]
  assign _T_54 = _T_51 ? _T_53 : _T_50; // @[LZD.scala 55:20]
  assign _T_55 = {_T_51,_T_54}; // @[Cat.scala 29:58]
  assign _T_56 = ~ _T_55; // @[convert.scala 21:22]
  assign _T_57 = realA[4:0]; // @[convert.scala 22:36]
  assign _T_58 = _T_56 < 3'h5; // @[Shift.scala 16:24]
  assign _T_60 = _T_56[2]; // @[Shift.scala 12:21]
  assign _T_61 = _T_57[0:0]; // @[Shift.scala 64:52]
  assign _T_63 = {_T_61,4'h0}; // @[Cat.scala 29:58]
  assign _T_64 = _T_60 ? _T_63 : _T_57; // @[Shift.scala 64:27]
  assign _T_65 = _T_56[1:0]; // @[Shift.scala 66:70]
  assign _T_66 = _T_65[1]; // @[Shift.scala 12:21]
  assign _T_67 = _T_64[2:0]; // @[Shift.scala 64:52]
  assign _T_69 = {_T_67,2'h0}; // @[Cat.scala 29:58]
  assign _T_70 = _T_66 ? _T_69 : _T_64; // @[Shift.scala 64:27]
  assign _T_71 = _T_65[0:0]; // @[Shift.scala 66:70]
  assign _T_73 = _T_70[3:0]; // @[Shift.scala 64:52]
  assign _T_74 = {_T_73,1'h0}; // @[Cat.scala 29:58]
  assign _T_75 = _T_71 ? _T_74 : _T_70; // @[Shift.scala 64:27]
  assign _T_76 = _T_58 ? _T_75 : 5'h0; // @[Shift.scala 16:10]
  assign _T_77 = _T_76[4:3]; // @[convert.scala 23:34]
  assign decA_fraction = _T_76[2:0]; // @[convert.scala 24:34]
  assign _T_79 = _T_15 == 1'h0; // @[convert.scala 25:26]
  assign _T_81 = _T_15 ? _T_56 : _T_55; // @[convert.scala 25:42]
  assign _T_84 = ~ _T_77; // @[convert.scala 26:67]
  assign _T_85 = _T_13 ? _T_84 : _T_77; // @[convert.scala 26:51]
  assign _T_86 = {_T_79,_T_81,_T_85}; // @[Cat.scala 29:58]
  assign _T_88 = realA[6:0]; // @[convert.scala 29:56]
  assign _T_89 = _T_88 != 7'h0; // @[convert.scala 29:60]
  assign _T_90 = ~ _T_89; // @[convert.scala 29:41]
  assign decA_isNaR = _T_13 & _T_90; // @[convert.scala 29:39]
  assign _T_93 = _T_13 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_93 & _T_90; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_86); // @[convert.scala 32:24]
  assign _T_102 = io_B[7]; // @[convert.scala 18:24]
  assign _T_103 = io_B[6]; // @[convert.scala 18:40]
  assign _T_104 = _T_102 ^ _T_103; // @[convert.scala 18:36]
  assign _T_105 = io_B[6:1]; // @[convert.scala 19:24]
  assign _T_106 = io_B[5:0]; // @[convert.scala 19:43]
  assign _T_107 = _T_105 ^ _T_106; // @[convert.scala 19:39]
  assign _T_108 = _T_107[5:2]; // @[LZD.scala 43:32]
  assign _T_109 = _T_108[3:2]; // @[LZD.scala 43:32]
  assign _T_110 = _T_109 != 2'h0; // @[LZD.scala 39:14]
  assign _T_111 = _T_109[1]; // @[LZD.scala 39:21]
  assign _T_112 = _T_109[0]; // @[LZD.scala 39:30]
  assign _T_113 = ~ _T_112; // @[LZD.scala 39:27]
  assign _T_114 = _T_111 | _T_113; // @[LZD.scala 39:25]
  assign _T_115 = {_T_110,_T_114}; // @[Cat.scala 29:58]
  assign _T_116 = _T_108[1:0]; // @[LZD.scala 44:32]
  assign _T_117 = _T_116 != 2'h0; // @[LZD.scala 39:14]
  assign _T_118 = _T_116[1]; // @[LZD.scala 39:21]
  assign _T_119 = _T_116[0]; // @[LZD.scala 39:30]
  assign _T_120 = ~ _T_119; // @[LZD.scala 39:27]
  assign _T_121 = _T_118 | _T_120; // @[LZD.scala 39:25]
  assign _T_122 = {_T_117,_T_121}; // @[Cat.scala 29:58]
  assign _T_123 = _T_115[1]; // @[Shift.scala 12:21]
  assign _T_124 = _T_122[1]; // @[Shift.scala 12:21]
  assign _T_125 = _T_123 | _T_124; // @[LZD.scala 49:16]
  assign _T_126 = ~ _T_124; // @[LZD.scala 49:27]
  assign _T_127 = _T_123 | _T_126; // @[LZD.scala 49:25]
  assign _T_128 = _T_115[0:0]; // @[LZD.scala 49:47]
  assign _T_129 = _T_122[0:0]; // @[LZD.scala 49:59]
  assign _T_130 = _T_123 ? _T_128 : _T_129; // @[LZD.scala 49:35]
  assign _T_132 = {_T_125,_T_127,_T_130}; // @[Cat.scala 29:58]
  assign _T_133 = _T_107[1:0]; // @[LZD.scala 44:32]
  assign _T_134 = _T_133 != 2'h0; // @[LZD.scala 39:14]
  assign _T_135 = _T_133[1]; // @[LZD.scala 39:21]
  assign _T_136 = _T_133[0]; // @[LZD.scala 39:30]
  assign _T_137 = ~ _T_136; // @[LZD.scala 39:27]
  assign _T_138 = _T_135 | _T_137; // @[LZD.scala 39:25]
  assign _T_139 = {_T_134,_T_138}; // @[Cat.scala 29:58]
  assign _T_140 = _T_132[2]; // @[Shift.scala 12:21]
  assign _T_142 = _T_132[1:0]; // @[LZD.scala 55:32]
  assign _T_143 = _T_140 ? _T_142 : _T_139; // @[LZD.scala 55:20]
  assign _T_144 = {_T_140,_T_143}; // @[Cat.scala 29:58]
  assign _T_145 = ~ _T_144; // @[convert.scala 21:22]
  assign _T_146 = io_B[4:0]; // @[convert.scala 22:36]
  assign _T_147 = _T_145 < 3'h5; // @[Shift.scala 16:24]
  assign _T_149 = _T_145[2]; // @[Shift.scala 12:21]
  assign _T_150 = _T_146[0:0]; // @[Shift.scala 64:52]
  assign _T_152 = {_T_150,4'h0}; // @[Cat.scala 29:58]
  assign _T_153 = _T_149 ? _T_152 : _T_146; // @[Shift.scala 64:27]
  assign _T_154 = _T_145[1:0]; // @[Shift.scala 66:70]
  assign _T_155 = _T_154[1]; // @[Shift.scala 12:21]
  assign _T_156 = _T_153[2:0]; // @[Shift.scala 64:52]
  assign _T_158 = {_T_156,2'h0}; // @[Cat.scala 29:58]
  assign _T_159 = _T_155 ? _T_158 : _T_153; // @[Shift.scala 64:27]
  assign _T_160 = _T_154[0:0]; // @[Shift.scala 66:70]
  assign _T_162 = _T_159[3:0]; // @[Shift.scala 64:52]
  assign _T_163 = {_T_162,1'h0}; // @[Cat.scala 29:58]
  assign _T_164 = _T_160 ? _T_163 : _T_159; // @[Shift.scala 64:27]
  assign _T_165 = _T_147 ? _T_164 : 5'h0; // @[Shift.scala 16:10]
  assign _T_166 = _T_165[4:3]; // @[convert.scala 23:34]
  assign decB_fraction = _T_165[2:0]; // @[convert.scala 24:34]
  assign _T_168 = _T_104 == 1'h0; // @[convert.scala 25:26]
  assign _T_170 = _T_104 ? _T_145 : _T_144; // @[convert.scala 25:42]
  assign _T_173 = ~ _T_166; // @[convert.scala 26:67]
  assign _T_174 = _T_102 ? _T_173 : _T_166; // @[convert.scala 26:51]
  assign _T_175 = {_T_168,_T_170,_T_174}; // @[Cat.scala 29:58]
  assign _T_177 = io_B[6:0]; // @[convert.scala 29:56]
  assign _T_178 = _T_177 != 7'h0; // @[convert.scala 29:60]
  assign _T_179 = ~ _T_178; // @[convert.scala 29:41]
  assign decB_isNaR = _T_102 & _T_179; // @[convert.scala 29:39]
  assign _T_182 = _T_102 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_182 & _T_179; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_175); // @[convert.scala 32:24]
  assign _T_191 = realC[7]; // @[convert.scala 18:24]
  assign _T_192 = realC[6]; // @[convert.scala 18:40]
  assign _T_193 = _T_191 ^ _T_192; // @[convert.scala 18:36]
  assign _T_194 = realC[6:1]; // @[convert.scala 19:24]
  assign _T_195 = realC[5:0]; // @[convert.scala 19:43]
  assign _T_196 = _T_194 ^ _T_195; // @[convert.scala 19:39]
  assign _T_197 = _T_196[5:2]; // @[LZD.scala 43:32]
  assign _T_198 = _T_197[3:2]; // @[LZD.scala 43:32]
  assign _T_199 = _T_198 != 2'h0; // @[LZD.scala 39:14]
  assign _T_200 = _T_198[1]; // @[LZD.scala 39:21]
  assign _T_201 = _T_198[0]; // @[LZD.scala 39:30]
  assign _T_202 = ~ _T_201; // @[LZD.scala 39:27]
  assign _T_203 = _T_200 | _T_202; // @[LZD.scala 39:25]
  assign _T_204 = {_T_199,_T_203}; // @[Cat.scala 29:58]
  assign _T_205 = _T_197[1:0]; // @[LZD.scala 44:32]
  assign _T_206 = _T_205 != 2'h0; // @[LZD.scala 39:14]
  assign _T_207 = _T_205[1]; // @[LZD.scala 39:21]
  assign _T_208 = _T_205[0]; // @[LZD.scala 39:30]
  assign _T_209 = ~ _T_208; // @[LZD.scala 39:27]
  assign _T_210 = _T_207 | _T_209; // @[LZD.scala 39:25]
  assign _T_211 = {_T_206,_T_210}; // @[Cat.scala 29:58]
  assign _T_212 = _T_204[1]; // @[Shift.scala 12:21]
  assign _T_213 = _T_211[1]; // @[Shift.scala 12:21]
  assign _T_214 = _T_212 | _T_213; // @[LZD.scala 49:16]
  assign _T_215 = ~ _T_213; // @[LZD.scala 49:27]
  assign _T_216 = _T_212 | _T_215; // @[LZD.scala 49:25]
  assign _T_217 = _T_204[0:0]; // @[LZD.scala 49:47]
  assign _T_218 = _T_211[0:0]; // @[LZD.scala 49:59]
  assign _T_219 = _T_212 ? _T_217 : _T_218; // @[LZD.scala 49:35]
  assign _T_221 = {_T_214,_T_216,_T_219}; // @[Cat.scala 29:58]
  assign _T_222 = _T_196[1:0]; // @[LZD.scala 44:32]
  assign _T_223 = _T_222 != 2'h0; // @[LZD.scala 39:14]
  assign _T_224 = _T_222[1]; // @[LZD.scala 39:21]
  assign _T_225 = _T_222[0]; // @[LZD.scala 39:30]
  assign _T_226 = ~ _T_225; // @[LZD.scala 39:27]
  assign _T_227 = _T_224 | _T_226; // @[LZD.scala 39:25]
  assign _T_228 = {_T_223,_T_227}; // @[Cat.scala 29:58]
  assign _T_229 = _T_221[2]; // @[Shift.scala 12:21]
  assign _T_231 = _T_221[1:0]; // @[LZD.scala 55:32]
  assign _T_232 = _T_229 ? _T_231 : _T_228; // @[LZD.scala 55:20]
  assign _T_233 = {_T_229,_T_232}; // @[Cat.scala 29:58]
  assign _T_234 = ~ _T_233; // @[convert.scala 21:22]
  assign _T_235 = realC[4:0]; // @[convert.scala 22:36]
  assign _T_236 = _T_234 < 3'h5; // @[Shift.scala 16:24]
  assign _T_238 = _T_234[2]; // @[Shift.scala 12:21]
  assign _T_239 = _T_235[0:0]; // @[Shift.scala 64:52]
  assign _T_241 = {_T_239,4'h0}; // @[Cat.scala 29:58]
  assign _T_242 = _T_238 ? _T_241 : _T_235; // @[Shift.scala 64:27]
  assign _T_243 = _T_234[1:0]; // @[Shift.scala 66:70]
  assign _T_244 = _T_243[1]; // @[Shift.scala 12:21]
  assign _T_245 = _T_242[2:0]; // @[Shift.scala 64:52]
  assign _T_247 = {_T_245,2'h0}; // @[Cat.scala 29:58]
  assign _T_248 = _T_244 ? _T_247 : _T_242; // @[Shift.scala 64:27]
  assign _T_249 = _T_243[0:0]; // @[Shift.scala 66:70]
  assign _T_251 = _T_248[3:0]; // @[Shift.scala 64:52]
  assign _T_252 = {_T_251,1'h0}; // @[Cat.scala 29:58]
  assign _T_253 = _T_249 ? _T_252 : _T_248; // @[Shift.scala 64:27]
  assign _T_254 = _T_236 ? _T_253 : 5'h0; // @[Shift.scala 16:10]
  assign _T_255 = _T_254[4:3]; // @[convert.scala 23:34]
  assign decC_fraction = _T_254[2:0]; // @[convert.scala 24:34]
  assign _T_257 = _T_193 == 1'h0; // @[convert.scala 25:26]
  assign _T_259 = _T_193 ? _T_234 : _T_233; // @[convert.scala 25:42]
  assign _T_262 = ~ _T_255; // @[convert.scala 26:67]
  assign _T_263 = _T_191 ? _T_262 : _T_255; // @[convert.scala 26:51]
  assign _T_264 = {_T_257,_T_259,_T_263}; // @[Cat.scala 29:58]
  assign _T_266 = realC[6:0]; // @[convert.scala 29:56]
  assign _T_267 = _T_266 != 7'h0; // @[convert.scala 29:60]
  assign _T_268 = ~ _T_267; // @[convert.scala 29:41]
  assign decC_isNaR = _T_191 & _T_268; // @[convert.scala 29:39]
  assign _T_271 = _T_191 == 1'h0; // @[convert.scala 30:19]
  assign decC_isZero = _T_271 & _T_268; // @[convert.scala 30:41]
  assign decC_scale = $signed(_T_264); // @[convert.scala 32:24]
  assign _T_279 = decA_isNaR | decB_isNaR; // @[PositFMA.scala 58:30]
  assign outIsNaR = _T_279 | decC_isNaR; // @[PositFMA.scala 58:44]
  assign _T_280 = ~ _T_13; // @[PositFMA.scala 59:34]
  assign _T_281 = ~ decA_isZero; // @[PositFMA.scala 59:47]
  assign _T_282 = _T_280 & _T_281; // @[PositFMA.scala 59:45]
  assign _T_284 = {_T_13,_T_282,decA_fraction}; // @[Cat.scala 29:58]
  assign sigA = $signed(_T_284); // @[PositFMA.scala 59:76]
  assign _T_285 = ~ _T_102; // @[PositFMA.scala 60:34]
  assign _T_286 = ~ decB_isZero; // @[PositFMA.scala 60:47]
  assign _T_287 = _T_285 & _T_286; // @[PositFMA.scala 60:45]
  assign _T_289 = {_T_102,_T_287,decB_fraction}; // @[Cat.scala 29:58]
  assign sigB = $signed(_T_289); // @[PositFMA.scala 60:76]
  assign _T_290 = $signed(sigA) * $signed(sigB); // @[PositFMA.scala 61:25]
  assign sigP = $unsigned(_T_290); // @[PositFMA.scala 61:33]
  assign head2 = sigP[9:8]; // @[PositFMA.scala 62:28]
  assign _T_291 = head2[1]; // @[PositFMA.scala 63:31]
  assign _T_292 = ~ _T_291; // @[PositFMA.scala 63:25]
  assign _T_293 = head2[0]; // @[PositFMA.scala 63:42]
  assign addTwo = _T_292 & _T_293; // @[PositFMA.scala 63:35]
  assign _T_294 = sigP[9]; // @[PositFMA.scala 65:23]
  assign _T_295 = sigP[7]; // @[PositFMA.scala 65:49]
  assign addOne = _T_294 ^ _T_295; // @[PositFMA.scala 65:43]
  assign _T_296 = {addTwo,addOne}; // @[Cat.scala 29:58]
  assign expBias = {1'b0,$signed(_T_296)}; // @[PositFMA.scala 66:39]
  assign mulSign = sigP[9:9]; // @[PositFMA.scala 67:28]
  assign _T_297 = $signed(decA_scale) + $signed(decB_scale); // @[PositFMA.scala 69:30]
  assign _GEN_12 = {{4{expBias[2]}},expBias}; // @[PositFMA.scala 69:44]
  assign _T_299 = $signed(_T_297) + $signed(_GEN_12); // @[PositFMA.scala 69:44]
  assign mulScale = $signed(_T_299); // @[PositFMA.scala 69:44]
  assign _T_300 = sigP[7:0]; // @[PositFMA.scala 72:29]
  assign _T_301 = sigP[6:0]; // @[PositFMA.scala 73:29]
  assign _T_302 = {_T_301, 1'h0}; // @[PositFMA.scala 73:48]
  assign mulSigTmp = addOne ? _T_300 : _T_302; // @[PositFMA.scala 70:22]
  assign _T_304 = mulSigTmp[7:7]; // @[PositFMA.scala 77:39]
  assign _T_305 = _T_304 | addTwo; // @[PositFMA.scala 77:43]
  assign _T_306 = mulSigTmp[6:0]; // @[PositFMA.scala 78:39]
  assign mulSig = {mulSign,_T_305,_T_306}; // @[Cat.scala 29:58]
  assign _T_332 = ~ addSign_phase2; // @[PositFMA.scala 107:29]
  assign _T_333 = ~ addZero_phase2; // @[PositFMA.scala 107:47]
  assign _T_334 = _T_332 & _T_333; // @[PositFMA.scala 107:45]
  assign extAddSig = {addSign_phase2,_T_334,addFrac_phase2,4'h0}; // @[Cat.scala 29:58]
  assign _GEN_13 = {{1{addScale_phase2[5]}},addScale_phase2}; // @[PositFMA.scala 111:39]
  assign mulGreater = $signed(mulScale_phase2) > $signed(_GEN_13); // @[PositFMA.scala 111:39]
  assign greaterScale = mulGreater ? $signed(mulScale_phase2) : $signed({{1{addScale_phase2[5]}},addScale_phase2}); // @[PositFMA.scala 112:26]
  assign smallerScale = mulGreater ? $signed({{1{addScale_phase2[5]}},addScale_phase2}) : $signed(mulScale_phase2); // @[PositFMA.scala 113:26]
  assign _T_338 = $signed(greaterScale) - $signed(smallerScale); // @[PositFMA.scala 114:36]
  assign scaleDiff = $signed(_T_338); // @[PositFMA.scala 114:36]
  assign greaterSig = mulGreater ? mulSig_phase2 : extAddSig; // @[PositFMA.scala 115:26]
  assign smallerSigTmp = mulGreater ? extAddSig : mulSig_phase2; // @[PositFMA.scala 116:26]
  assign _T_339 = $unsigned(scaleDiff); // @[PositFMA.scala 117:69]
  assign _T_340 = _T_339 < 7'h9; // @[Shift.scala 39:24]
  assign _T_341 = _T_339[3:0]; // @[Shift.scala 40:44]
  assign _T_342 = smallerSigTmp[8:8]; // @[Shift.scala 90:30]
  assign _T_343 = smallerSigTmp[7:0]; // @[Shift.scala 90:48]
  assign _T_344 = _T_343 != 8'h0; // @[Shift.scala 90:57]
  assign _T_345 = _T_342 | _T_344; // @[Shift.scala 90:39]
  assign _T_346 = _T_341[3]; // @[Shift.scala 12:21]
  assign _T_347 = smallerSigTmp[8]; // @[Shift.scala 12:21]
  assign _T_349 = _T_347 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_350 = {_T_349,_T_345}; // @[Cat.scala 29:58]
  assign _T_351 = _T_346 ? _T_350 : smallerSigTmp; // @[Shift.scala 91:22]
  assign _T_352 = _T_341[2:0]; // @[Shift.scala 92:77]
  assign _T_353 = _T_351[8:4]; // @[Shift.scala 90:30]
  assign _T_354 = _T_351[3:0]; // @[Shift.scala 90:48]
  assign _T_355 = _T_354 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_14 = {{4'd0}, _T_355}; // @[Shift.scala 90:39]
  assign _T_356 = _T_353 | _GEN_14; // @[Shift.scala 90:39]
  assign _T_357 = _T_352[2]; // @[Shift.scala 12:21]
  assign _T_358 = _T_351[8]; // @[Shift.scala 12:21]
  assign _T_360 = _T_358 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_361 = {_T_360,_T_356}; // @[Cat.scala 29:58]
  assign _T_362 = _T_357 ? _T_361 : _T_351; // @[Shift.scala 91:22]
  assign _T_363 = _T_352[1:0]; // @[Shift.scala 92:77]
  assign _T_364 = _T_362[8:2]; // @[Shift.scala 90:30]
  assign _T_365 = _T_362[1:0]; // @[Shift.scala 90:48]
  assign _T_366 = _T_365 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_15 = {{6'd0}, _T_366}; // @[Shift.scala 90:39]
  assign _T_367 = _T_364 | _GEN_15; // @[Shift.scala 90:39]
  assign _T_368 = _T_363[1]; // @[Shift.scala 12:21]
  assign _T_369 = _T_362[8]; // @[Shift.scala 12:21]
  assign _T_371 = _T_369 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_372 = {_T_371,_T_367}; // @[Cat.scala 29:58]
  assign _T_373 = _T_368 ? _T_372 : _T_362; // @[Shift.scala 91:22]
  assign _T_374 = _T_363[0:0]; // @[Shift.scala 92:77]
  assign _T_375 = _T_373[8:1]; // @[Shift.scala 90:30]
  assign _T_376 = _T_373[0:0]; // @[Shift.scala 90:48]
  assign _GEN_16 = {{7'd0}, _T_376}; // @[Shift.scala 90:39]
  assign _T_378 = _T_375 | _GEN_16; // @[Shift.scala 90:39]
  assign _T_380 = _T_373[8]; // @[Shift.scala 12:21]
  assign _T_381 = {_T_380,_T_378}; // @[Cat.scala 29:58]
  assign _T_382 = _T_374 ? _T_381 : _T_373; // @[Shift.scala 91:22]
  assign _T_385 = _T_347 ? 9'h1ff : 9'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_340 ? _T_382 : _T_385; // @[Shift.scala 39:10]
  assign rawSumSig = greaterSig + smallerSig; // @[PositFMA.scala 118:34]
  assign _T_386 = mulSig_phase2[8:8]; // @[PositFMA.scala 119:42]
  assign _T_387 = _T_386 ^ addSign_phase2; // @[PositFMA.scala 119:46]
  assign _T_388 = rawSumSig[9:9]; // @[PositFMA.scala 119:79]
  assign sumSign = _T_387 ^ _T_388; // @[PositFMA.scala 119:63]
  assign _T_390 = greaterSig + smallerSig; // @[PositFMA.scala 120:50]
  assign signSumSig = {sumSign,_T_390}; // @[Cat.scala 29:58]
  assign _T_391 = signSumSig[9:1]; // @[PositFMA.scala 124:33]
  assign _T_392 = signSumSig[8:0]; // @[PositFMA.scala 124:68]
  assign sumXor = _T_391 ^ _T_392; // @[PositFMA.scala 124:51]
  assign _T_393 = sumXor[8:1]; // @[LZD.scala 43:32]
  assign _T_394 = _T_393[7:4]; // @[LZD.scala 43:32]
  assign _T_395 = _T_394[3:2]; // @[LZD.scala 43:32]
  assign _T_396 = _T_395 != 2'h0; // @[LZD.scala 39:14]
  assign _T_397 = _T_395[1]; // @[LZD.scala 39:21]
  assign _T_398 = _T_395[0]; // @[LZD.scala 39:30]
  assign _T_399 = ~ _T_398; // @[LZD.scala 39:27]
  assign _T_400 = _T_397 | _T_399; // @[LZD.scala 39:25]
  assign _T_401 = {_T_396,_T_400}; // @[Cat.scala 29:58]
  assign _T_402 = _T_394[1:0]; // @[LZD.scala 44:32]
  assign _T_403 = _T_402 != 2'h0; // @[LZD.scala 39:14]
  assign _T_404 = _T_402[1]; // @[LZD.scala 39:21]
  assign _T_405 = _T_402[0]; // @[LZD.scala 39:30]
  assign _T_406 = ~ _T_405; // @[LZD.scala 39:27]
  assign _T_407 = _T_404 | _T_406; // @[LZD.scala 39:25]
  assign _T_408 = {_T_403,_T_407}; // @[Cat.scala 29:58]
  assign _T_409 = _T_401[1]; // @[Shift.scala 12:21]
  assign _T_410 = _T_408[1]; // @[Shift.scala 12:21]
  assign _T_411 = _T_409 | _T_410; // @[LZD.scala 49:16]
  assign _T_412 = ~ _T_410; // @[LZD.scala 49:27]
  assign _T_413 = _T_409 | _T_412; // @[LZD.scala 49:25]
  assign _T_414 = _T_401[0:0]; // @[LZD.scala 49:47]
  assign _T_415 = _T_408[0:0]; // @[LZD.scala 49:59]
  assign _T_416 = _T_409 ? _T_414 : _T_415; // @[LZD.scala 49:35]
  assign _T_418 = {_T_411,_T_413,_T_416}; // @[Cat.scala 29:58]
  assign _T_419 = _T_393[3:0]; // @[LZD.scala 44:32]
  assign _T_420 = _T_419[3:2]; // @[LZD.scala 43:32]
  assign _T_421 = _T_420 != 2'h0; // @[LZD.scala 39:14]
  assign _T_422 = _T_420[1]; // @[LZD.scala 39:21]
  assign _T_423 = _T_420[0]; // @[LZD.scala 39:30]
  assign _T_424 = ~ _T_423; // @[LZD.scala 39:27]
  assign _T_425 = _T_422 | _T_424; // @[LZD.scala 39:25]
  assign _T_426 = {_T_421,_T_425}; // @[Cat.scala 29:58]
  assign _T_427 = _T_419[1:0]; // @[LZD.scala 44:32]
  assign _T_428 = _T_427 != 2'h0; // @[LZD.scala 39:14]
  assign _T_429 = _T_427[1]; // @[LZD.scala 39:21]
  assign _T_430 = _T_427[0]; // @[LZD.scala 39:30]
  assign _T_431 = ~ _T_430; // @[LZD.scala 39:27]
  assign _T_432 = _T_429 | _T_431; // @[LZD.scala 39:25]
  assign _T_433 = {_T_428,_T_432}; // @[Cat.scala 29:58]
  assign _T_434 = _T_426[1]; // @[Shift.scala 12:21]
  assign _T_435 = _T_433[1]; // @[Shift.scala 12:21]
  assign _T_436 = _T_434 | _T_435; // @[LZD.scala 49:16]
  assign _T_437 = ~ _T_435; // @[LZD.scala 49:27]
  assign _T_438 = _T_434 | _T_437; // @[LZD.scala 49:25]
  assign _T_439 = _T_426[0:0]; // @[LZD.scala 49:47]
  assign _T_440 = _T_433[0:0]; // @[LZD.scala 49:59]
  assign _T_441 = _T_434 ? _T_439 : _T_440; // @[LZD.scala 49:35]
  assign _T_443 = {_T_436,_T_438,_T_441}; // @[Cat.scala 29:58]
  assign _T_444 = _T_418[2]; // @[Shift.scala 12:21]
  assign _T_445 = _T_443[2]; // @[Shift.scala 12:21]
  assign _T_446 = _T_444 | _T_445; // @[LZD.scala 49:16]
  assign _T_447 = ~ _T_445; // @[LZD.scala 49:27]
  assign _T_448 = _T_444 | _T_447; // @[LZD.scala 49:25]
  assign _T_449 = _T_418[1:0]; // @[LZD.scala 49:47]
  assign _T_450 = _T_443[1:0]; // @[LZD.scala 49:59]
  assign _T_451 = _T_444 ? _T_449 : _T_450; // @[LZD.scala 49:35]
  assign _T_453 = {_T_446,_T_448,_T_451}; // @[Cat.scala 29:58]
  assign _T_454 = sumXor[0:0]; // @[LZD.scala 44:32]
  assign _T_456 = _T_453[3]; // @[Shift.scala 12:21]
  assign _T_459 = {2'h3,_T_454}; // @[Cat.scala 29:58]
  assign _T_460 = _T_453[2:0]; // @[LZD.scala 55:32]
  assign _T_461 = _T_456 ? _T_460 : _T_459; // @[LZD.scala 55:20]
  assign sumLZD = {_T_456,_T_461}; // @[Cat.scala 29:58]
  assign shiftValue = ~ sumLZD; // @[PositFMA.scala 126:24]
  assign _T_462 = signSumSig[7:0]; // @[PositFMA.scala 127:38]
  assign _T_463 = shiftValue < 4'h8; // @[Shift.scala 16:24]
  assign _T_464 = shiftValue[2:0]; // @[Shift.scala 17:37]
  assign _T_465 = _T_464[2]; // @[Shift.scala 12:21]
  assign _T_466 = _T_462[3:0]; // @[Shift.scala 64:52]
  assign _T_468 = {_T_466,4'h0}; // @[Cat.scala 29:58]
  assign _T_469 = _T_465 ? _T_468 : _T_462; // @[Shift.scala 64:27]
  assign _T_470 = _T_464[1:0]; // @[Shift.scala 66:70]
  assign _T_471 = _T_470[1]; // @[Shift.scala 12:21]
  assign _T_472 = _T_469[5:0]; // @[Shift.scala 64:52]
  assign _T_474 = {_T_472,2'h0}; // @[Cat.scala 29:58]
  assign _T_475 = _T_471 ? _T_474 : _T_469; // @[Shift.scala 64:27]
  assign _T_476 = _T_470[0:0]; // @[Shift.scala 66:70]
  assign _T_478 = _T_475[6:0]; // @[Shift.scala 64:52]
  assign _T_479 = {_T_478,1'h0}; // @[Cat.scala 29:58]
  assign _T_480 = _T_476 ? _T_479 : _T_475; // @[Shift.scala 64:27]
  assign normalFracTmp = _T_463 ? _T_480 : 8'h0; // @[Shift.scala 16:10]
  assign _T_482 = $signed(greaterScale) + $signed(7'sh2); // @[PositFMA.scala 130:36]
  assign _T_483 = $signed(_T_482); // @[PositFMA.scala 130:36]
  assign _T_484 = {1'h1,_T_456,_T_461}; // @[Cat.scala 29:58]
  assign _T_485 = $signed(_T_484); // @[PositFMA.scala 130:61]
  assign _GEN_17 = {{2{_T_485[4]}},_T_485}; // @[PositFMA.scala 130:42]
  assign _T_487 = $signed(_T_483) + $signed(_GEN_17); // @[PositFMA.scala 130:42]
  assign sumScale = $signed(_T_487); // @[PositFMA.scala 130:42]
  assign sumFrac = normalFracTmp[7:5]; // @[PositFMA.scala 131:41]
  assign grsTmp = normalFracTmp[4:0]; // @[PositFMA.scala 134:41]
  assign _T_488 = grsTmp[4:3]; // @[PositFMA.scala 137:40]
  assign _T_489 = grsTmp[2:0]; // @[PositFMA.scala 137:56]
  assign _T_490 = _T_489 != 3'h0; // @[PositFMA.scala 137:60]
  assign underflow = $signed(sumScale) < $signed(-7'sh19); // @[PositFMA.scala 144:32]
  assign overflow = $signed(sumScale) > $signed(7'sh18); // @[PositFMA.scala 145:32]
  assign _T_491 = signSumSig != 10'h0; // @[PositFMA.scala 154:32]
  assign decF_isZero = ~ _T_491; // @[PositFMA.scala 154:20]
  assign _T_493 = underflow ? $signed(-7'sh19) : $signed(sumScale); // @[Mux.scala 87:16]
  assign _T_494 = overflow ? $signed(7'sh18) : $signed(_T_493); // @[Mux.scala 87:16]
  assign _GEN_18 = _T_494[5:0]; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  assign decF_scale = $signed(_GEN_18); // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  assign _T_495 = decF_scale[1:0]; // @[convert.scala 46:61]
  assign _T_496 = ~ _T_495; // @[convert.scala 46:52]
  assign _T_498 = sumSign ? _T_496 : _T_495; // @[convert.scala 46:42]
  assign _T_499 = decF_scale[5:2]; // @[convert.scala 48:34]
  assign _T_500 = _T_499[3:3]; // @[convert.scala 49:36]
  assign _T_502 = ~ _T_499; // @[convert.scala 50:36]
  assign _T_503 = $signed(_T_502); // @[convert.scala 50:36]
  assign _T_504 = _T_500 ? $signed(_T_503) : $signed(_T_499); // @[convert.scala 50:28]
  assign _T_505 = _T_500 ^ sumSign; // @[convert.scala 51:31]
  assign _T_506 = ~ _T_505; // @[convert.scala 52:43]
  assign _T_510 = {_T_506,_T_505,_T_498,sumFrac,_T_488,_T_490}; // @[Cat.scala 29:58]
  assign _T_511 = $unsigned(_T_504); // @[Shift.scala 39:17]
  assign _T_512 = _T_511 < 4'ha; // @[Shift.scala 39:24]
  assign _T_514 = _T_510[9:8]; // @[Shift.scala 90:30]
  assign _T_515 = _T_510[7:0]; // @[Shift.scala 90:48]
  assign _T_516 = _T_515 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_19 = {{1'd0}, _T_516}; // @[Shift.scala 90:39]
  assign _T_517 = _T_514 | _GEN_19; // @[Shift.scala 90:39]
  assign _T_518 = _T_511[3]; // @[Shift.scala 12:21]
  assign _T_519 = _T_510[9]; // @[Shift.scala 12:21]
  assign _T_521 = _T_519 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_522 = {_T_521,_T_517}; // @[Cat.scala 29:58]
  assign _T_523 = _T_518 ? _T_522 : _T_510; // @[Shift.scala 91:22]
  assign _T_524 = _T_511[2:0]; // @[Shift.scala 92:77]
  assign _T_525 = _T_523[9:4]; // @[Shift.scala 90:30]
  assign _T_526 = _T_523[3:0]; // @[Shift.scala 90:48]
  assign _T_527 = _T_526 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_20 = {{5'd0}, _T_527}; // @[Shift.scala 90:39]
  assign _T_528 = _T_525 | _GEN_20; // @[Shift.scala 90:39]
  assign _T_529 = _T_524[2]; // @[Shift.scala 12:21]
  assign _T_530 = _T_523[9]; // @[Shift.scala 12:21]
  assign _T_532 = _T_530 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_533 = {_T_532,_T_528}; // @[Cat.scala 29:58]
  assign _T_534 = _T_529 ? _T_533 : _T_523; // @[Shift.scala 91:22]
  assign _T_535 = _T_524[1:0]; // @[Shift.scala 92:77]
  assign _T_536 = _T_534[9:2]; // @[Shift.scala 90:30]
  assign _T_537 = _T_534[1:0]; // @[Shift.scala 90:48]
  assign _T_538 = _T_537 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_21 = {{7'd0}, _T_538}; // @[Shift.scala 90:39]
  assign _T_539 = _T_536 | _GEN_21; // @[Shift.scala 90:39]
  assign _T_540 = _T_535[1]; // @[Shift.scala 12:21]
  assign _T_541 = _T_534[9]; // @[Shift.scala 12:21]
  assign _T_543 = _T_541 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_544 = {_T_543,_T_539}; // @[Cat.scala 29:58]
  assign _T_545 = _T_540 ? _T_544 : _T_534; // @[Shift.scala 91:22]
  assign _T_546 = _T_535[0:0]; // @[Shift.scala 92:77]
  assign _T_547 = _T_545[9:1]; // @[Shift.scala 90:30]
  assign _T_548 = _T_545[0:0]; // @[Shift.scala 90:48]
  assign _GEN_22 = {{8'd0}, _T_548}; // @[Shift.scala 90:39]
  assign _T_550 = _T_547 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_552 = _T_545[9]; // @[Shift.scala 12:21]
  assign _T_553 = {_T_552,_T_550}; // @[Cat.scala 29:58]
  assign _T_554 = _T_546 ? _T_553 : _T_545; // @[Shift.scala 91:22]
  assign _T_557 = _T_519 ? 10'h3ff : 10'h0; // @[Bitwise.scala 71:12]
  assign _T_558 = _T_512 ? _T_554 : _T_557; // @[Shift.scala 39:10]
  assign _T_559 = _T_558[3]; // @[convert.scala 55:31]
  assign _T_560 = _T_558[2]; // @[convert.scala 56:31]
  assign _T_561 = _T_558[1]; // @[convert.scala 57:31]
  assign _T_562 = _T_558[0]; // @[convert.scala 58:31]
  assign _T_563 = _T_558[9:3]; // @[convert.scala 59:69]
  assign _T_564 = _T_563 != 7'h0; // @[convert.scala 59:81]
  assign _T_565 = ~ _T_564; // @[convert.scala 59:50]
  assign _T_567 = _T_563 == 7'h7f; // @[convert.scala 60:81]
  assign _T_568 = _T_559 | _T_561; // @[convert.scala 61:44]
  assign _T_569 = _T_568 | _T_562; // @[convert.scala 61:52]
  assign _T_570 = _T_560 & _T_569; // @[convert.scala 61:36]
  assign _T_571 = ~ _T_567; // @[convert.scala 62:63]
  assign _T_572 = _T_571 & _T_570; // @[convert.scala 62:103]
  assign _T_573 = _T_565 | _T_572; // @[convert.scala 62:60]
  assign _GEN_23 = {{6'd0}, _T_573}; // @[convert.scala 63:56]
  assign _T_576 = _T_563 + _GEN_23; // @[convert.scala 63:56]
  assign _T_577 = {sumSign,_T_576}; // @[Cat.scala 29:58]
  assign io_F = _T_585; // @[PositFMA.scala 174:15]
  assign io_outValid = _T_581; // @[PositFMA.scala 173:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  outIsNaR_phase2 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mulSig_phase2 = _RAND_1[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  addFrac_phase2 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mulScale_phase2 = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addScale_phase2 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addSign_phase2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addZero_phase2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  inValid_phase2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_581 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_585 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (io_inValid) begin
      outIsNaR_phase2 <= outIsNaR;
    end
    if (io_inValid) begin
      mulSig_phase2 <= mulSig;
    end
    if (io_inValid) begin
      addFrac_phase2 <= decC_fraction;
    end
    if (io_inValid) begin
      mulScale_phase2 <= mulScale;
    end
    if (io_inValid) begin
      addScale_phase2 <= decC_scale;
    end
    if (io_inValid) begin
      addSign_phase2 <= _T_191;
    end
    if (io_inValid) begin
      addZero_phase2 <= decC_isZero;
    end
    if (reset) begin
      inValid_phase2 <= 1'h0;
    end else begin
      inValid_phase2 <= io_inValid;
    end
    if (reset) begin
      _T_581 <= 1'h0;
    end else begin
      _T_581 <= inValid_phase2;
    end
    if (inValid_phase2) begin
      if (outIsNaR_phase2) begin
        _T_585 <= 8'h80;
      end else begin
        if (decF_isZero) begin
          _T_585 <= 8'h0;
        end else begin
          _T_585 <= _T_577;
        end
      end
    end
  end
endmodule
