module PositFMA14_1(
  input         clock,
  input         reset,
  input         io_inValid,
  input  [1:0]  io_fmaOp,
  input  [13:0] io_A,
  input  [13:0] io_B,
  input  [13:0] io_C,
  output [13:0] io_F,
  output        io_outValid
);
  wire  _T; // @[PositFMA.scala 47:36]
  wire [13:0] _T_2; // @[Bitwise.scala 71:12]
  wire [13:0] _T_3; // @[PositFMA.scala 47:41]
  wire [13:0] _GEN_10; // @[PositFMA.scala 47:49]
  wire [13:0] realA; // @[PositFMA.scala 47:49]
  wire  _T_6; // @[PositFMA.scala 48:36]
  wire [13:0] _T_8; // @[Bitwise.scala 71:12]
  wire [13:0] _T_9; // @[PositFMA.scala 48:41]
  wire [13:0] _GEN_11; // @[PositFMA.scala 48:49]
  wire [13:0] realC; // @[PositFMA.scala 48:49]
  wire  _T_13; // @[convert.scala 18:24]
  wire  _T_14; // @[convert.scala 18:40]
  wire  _T_15; // @[convert.scala 18:36]
  wire [11:0] _T_16; // @[convert.scala 19:24]
  wire [11:0] _T_17; // @[convert.scala 19:43]
  wire [11:0] _T_18; // @[convert.scala 19:39]
  wire [7:0] _T_19; // @[LZD.scala 43:32]
  wire [3:0] _T_20; // @[LZD.scala 43:32]
  wire [1:0] _T_21; // @[LZD.scala 43:32]
  wire  _T_22; // @[LZD.scala 39:14]
  wire  _T_23; // @[LZD.scala 39:21]
  wire  _T_24; // @[LZD.scala 39:30]
  wire  _T_25; // @[LZD.scala 39:27]
  wire  _T_26; // @[LZD.scala 39:25]
  wire [1:0] _T_27; // @[Cat.scala 29:58]
  wire [1:0] _T_28; // @[LZD.scala 44:32]
  wire  _T_29; // @[LZD.scala 39:14]
  wire  _T_30; // @[LZD.scala 39:21]
  wire  _T_31; // @[LZD.scala 39:30]
  wire  _T_32; // @[LZD.scala 39:27]
  wire  _T_33; // @[LZD.scala 39:25]
  wire [1:0] _T_34; // @[Cat.scala 29:58]
  wire  _T_35; // @[Shift.scala 12:21]
  wire  _T_36; // @[Shift.scala 12:21]
  wire  _T_37; // @[LZD.scala 49:16]
  wire  _T_38; // @[LZD.scala 49:27]
  wire  _T_39; // @[LZD.scala 49:25]
  wire  _T_40; // @[LZD.scala 49:47]
  wire  _T_41; // @[LZD.scala 49:59]
  wire  _T_42; // @[LZD.scala 49:35]
  wire [2:0] _T_44; // @[Cat.scala 29:58]
  wire [3:0] _T_45; // @[LZD.scala 44:32]
  wire [1:0] _T_46; // @[LZD.scala 43:32]
  wire  _T_47; // @[LZD.scala 39:14]
  wire  _T_48; // @[LZD.scala 39:21]
  wire  _T_49; // @[LZD.scala 39:30]
  wire  _T_50; // @[LZD.scala 39:27]
  wire  _T_51; // @[LZD.scala 39:25]
  wire [1:0] _T_52; // @[Cat.scala 29:58]
  wire [1:0] _T_53; // @[LZD.scala 44:32]
  wire  _T_54; // @[LZD.scala 39:14]
  wire  _T_55; // @[LZD.scala 39:21]
  wire  _T_56; // @[LZD.scala 39:30]
  wire  _T_57; // @[LZD.scala 39:27]
  wire  _T_58; // @[LZD.scala 39:25]
  wire [1:0] _T_59; // @[Cat.scala 29:58]
  wire  _T_60; // @[Shift.scala 12:21]
  wire  _T_61; // @[Shift.scala 12:21]
  wire  _T_62; // @[LZD.scala 49:16]
  wire  _T_63; // @[LZD.scala 49:27]
  wire  _T_64; // @[LZD.scala 49:25]
  wire  _T_65; // @[LZD.scala 49:47]
  wire  _T_66; // @[LZD.scala 49:59]
  wire  _T_67; // @[LZD.scala 49:35]
  wire [2:0] _T_69; // @[Cat.scala 29:58]
  wire  _T_70; // @[Shift.scala 12:21]
  wire  _T_71; // @[Shift.scala 12:21]
  wire  _T_72; // @[LZD.scala 49:16]
  wire  _T_73; // @[LZD.scala 49:27]
  wire  _T_74; // @[LZD.scala 49:25]
  wire [1:0] _T_75; // @[LZD.scala 49:47]
  wire [1:0] _T_76; // @[LZD.scala 49:59]
  wire [1:0] _T_77; // @[LZD.scala 49:35]
  wire [3:0] _T_79; // @[Cat.scala 29:58]
  wire [3:0] _T_80; // @[LZD.scala 44:32]
  wire [1:0] _T_81; // @[LZD.scala 43:32]
  wire  _T_82; // @[LZD.scala 39:14]
  wire  _T_83; // @[LZD.scala 39:21]
  wire  _T_84; // @[LZD.scala 39:30]
  wire  _T_85; // @[LZD.scala 39:27]
  wire  _T_86; // @[LZD.scala 39:25]
  wire [1:0] _T_87; // @[Cat.scala 29:58]
  wire [1:0] _T_88; // @[LZD.scala 44:32]
  wire  _T_89; // @[LZD.scala 39:14]
  wire  _T_90; // @[LZD.scala 39:21]
  wire  _T_91; // @[LZD.scala 39:30]
  wire  _T_92; // @[LZD.scala 39:27]
  wire  _T_93; // @[LZD.scala 39:25]
  wire [1:0] _T_94; // @[Cat.scala 29:58]
  wire  _T_95; // @[Shift.scala 12:21]
  wire  _T_96; // @[Shift.scala 12:21]
  wire  _T_97; // @[LZD.scala 49:16]
  wire  _T_98; // @[LZD.scala 49:27]
  wire  _T_99; // @[LZD.scala 49:25]
  wire  _T_100; // @[LZD.scala 49:47]
  wire  _T_101; // @[LZD.scala 49:59]
  wire  _T_102; // @[LZD.scala 49:35]
  wire [2:0] _T_104; // @[Cat.scala 29:58]
  wire  _T_105; // @[Shift.scala 12:21]
  wire [2:0] _T_107; // @[LZD.scala 55:32]
  wire [2:0] _T_108; // @[LZD.scala 55:20]
  wire [3:0] _T_109; // @[Cat.scala 29:58]
  wire [3:0] _T_110; // @[convert.scala 21:22]
  wire [10:0] _T_111; // @[convert.scala 22:36]
  wire  _T_112; // @[Shift.scala 16:24]
  wire  _T_114; // @[Shift.scala 12:21]
  wire [2:0] _T_115; // @[Shift.scala 64:52]
  wire [10:0] _T_117; // @[Cat.scala 29:58]
  wire [10:0] _T_118; // @[Shift.scala 64:27]
  wire [2:0] _T_119; // @[Shift.scala 66:70]
  wire  _T_120; // @[Shift.scala 12:21]
  wire [6:0] _T_121; // @[Shift.scala 64:52]
  wire [10:0] _T_123; // @[Cat.scala 29:58]
  wire [10:0] _T_124; // @[Shift.scala 64:27]
  wire [1:0] _T_125; // @[Shift.scala 66:70]
  wire  _T_126; // @[Shift.scala 12:21]
  wire [8:0] _T_127; // @[Shift.scala 64:52]
  wire [10:0] _T_129; // @[Cat.scala 29:58]
  wire [10:0] _T_130; // @[Shift.scala 64:27]
  wire  _T_131; // @[Shift.scala 66:70]
  wire [9:0] _T_133; // @[Shift.scala 64:52]
  wire [10:0] _T_134; // @[Cat.scala 29:58]
  wire [10:0] _T_135; // @[Shift.scala 64:27]
  wire [10:0] _T_136; // @[Shift.scala 16:10]
  wire  _T_137; // @[convert.scala 23:34]
  wire [9:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_139; // @[convert.scala 25:26]
  wire [3:0] _T_141; // @[convert.scala 25:42]
  wire  _T_144; // @[convert.scala 26:67]
  wire  _T_145; // @[convert.scala 26:51]
  wire [5:0] _T_146; // @[Cat.scala 29:58]
  wire [12:0] _T_148; // @[convert.scala 29:56]
  wire  _T_149; // @[convert.scala 29:60]
  wire  _T_150; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_153; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [5:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_162; // @[convert.scala 18:24]
  wire  _T_163; // @[convert.scala 18:40]
  wire  _T_164; // @[convert.scala 18:36]
  wire [11:0] _T_165; // @[convert.scala 19:24]
  wire [11:0] _T_166; // @[convert.scala 19:43]
  wire [11:0] _T_167; // @[convert.scala 19:39]
  wire [7:0] _T_168; // @[LZD.scala 43:32]
  wire [3:0] _T_169; // @[LZD.scala 43:32]
  wire [1:0] _T_170; // @[LZD.scala 43:32]
  wire  _T_171; // @[LZD.scala 39:14]
  wire  _T_172; // @[LZD.scala 39:21]
  wire  _T_173; // @[LZD.scala 39:30]
  wire  _T_174; // @[LZD.scala 39:27]
  wire  _T_175; // @[LZD.scala 39:25]
  wire [1:0] _T_176; // @[Cat.scala 29:58]
  wire [1:0] _T_177; // @[LZD.scala 44:32]
  wire  _T_178; // @[LZD.scala 39:14]
  wire  _T_179; // @[LZD.scala 39:21]
  wire  _T_180; // @[LZD.scala 39:30]
  wire  _T_181; // @[LZD.scala 39:27]
  wire  _T_182; // @[LZD.scala 39:25]
  wire [1:0] _T_183; // @[Cat.scala 29:58]
  wire  _T_184; // @[Shift.scala 12:21]
  wire  _T_185; // @[Shift.scala 12:21]
  wire  _T_186; // @[LZD.scala 49:16]
  wire  _T_187; // @[LZD.scala 49:27]
  wire  _T_188; // @[LZD.scala 49:25]
  wire  _T_189; // @[LZD.scala 49:47]
  wire  _T_190; // @[LZD.scala 49:59]
  wire  _T_191; // @[LZD.scala 49:35]
  wire [2:0] _T_193; // @[Cat.scala 29:58]
  wire [3:0] _T_194; // @[LZD.scala 44:32]
  wire [1:0] _T_195; // @[LZD.scala 43:32]
  wire  _T_196; // @[LZD.scala 39:14]
  wire  _T_197; // @[LZD.scala 39:21]
  wire  _T_198; // @[LZD.scala 39:30]
  wire  _T_199; // @[LZD.scala 39:27]
  wire  _T_200; // @[LZD.scala 39:25]
  wire [1:0] _T_201; // @[Cat.scala 29:58]
  wire [1:0] _T_202; // @[LZD.scala 44:32]
  wire  _T_203; // @[LZD.scala 39:14]
  wire  _T_204; // @[LZD.scala 39:21]
  wire  _T_205; // @[LZD.scala 39:30]
  wire  _T_206; // @[LZD.scala 39:27]
  wire  _T_207; // @[LZD.scala 39:25]
  wire [1:0] _T_208; // @[Cat.scala 29:58]
  wire  _T_209; // @[Shift.scala 12:21]
  wire  _T_210; // @[Shift.scala 12:21]
  wire  _T_211; // @[LZD.scala 49:16]
  wire  _T_212; // @[LZD.scala 49:27]
  wire  _T_213; // @[LZD.scala 49:25]
  wire  _T_214; // @[LZD.scala 49:47]
  wire  _T_215; // @[LZD.scala 49:59]
  wire  _T_216; // @[LZD.scala 49:35]
  wire [2:0] _T_218; // @[Cat.scala 29:58]
  wire  _T_219; // @[Shift.scala 12:21]
  wire  _T_220; // @[Shift.scala 12:21]
  wire  _T_221; // @[LZD.scala 49:16]
  wire  _T_222; // @[LZD.scala 49:27]
  wire  _T_223; // @[LZD.scala 49:25]
  wire [1:0] _T_224; // @[LZD.scala 49:47]
  wire [1:0] _T_225; // @[LZD.scala 49:59]
  wire [1:0] _T_226; // @[LZD.scala 49:35]
  wire [3:0] _T_228; // @[Cat.scala 29:58]
  wire [3:0] _T_229; // @[LZD.scala 44:32]
  wire [1:0] _T_230; // @[LZD.scala 43:32]
  wire  _T_231; // @[LZD.scala 39:14]
  wire  _T_232; // @[LZD.scala 39:21]
  wire  _T_233; // @[LZD.scala 39:30]
  wire  _T_234; // @[LZD.scala 39:27]
  wire  _T_235; // @[LZD.scala 39:25]
  wire [1:0] _T_236; // @[Cat.scala 29:58]
  wire [1:0] _T_237; // @[LZD.scala 44:32]
  wire  _T_238; // @[LZD.scala 39:14]
  wire  _T_239; // @[LZD.scala 39:21]
  wire  _T_240; // @[LZD.scala 39:30]
  wire  _T_241; // @[LZD.scala 39:27]
  wire  _T_242; // @[LZD.scala 39:25]
  wire [1:0] _T_243; // @[Cat.scala 29:58]
  wire  _T_244; // @[Shift.scala 12:21]
  wire  _T_245; // @[Shift.scala 12:21]
  wire  _T_246; // @[LZD.scala 49:16]
  wire  _T_247; // @[LZD.scala 49:27]
  wire  _T_248; // @[LZD.scala 49:25]
  wire  _T_249; // @[LZD.scala 49:47]
  wire  _T_250; // @[LZD.scala 49:59]
  wire  _T_251; // @[LZD.scala 49:35]
  wire [2:0] _T_253; // @[Cat.scala 29:58]
  wire  _T_254; // @[Shift.scala 12:21]
  wire [2:0] _T_256; // @[LZD.scala 55:32]
  wire [2:0] _T_257; // @[LZD.scala 55:20]
  wire [3:0] _T_258; // @[Cat.scala 29:58]
  wire [3:0] _T_259; // @[convert.scala 21:22]
  wire [10:0] _T_260; // @[convert.scala 22:36]
  wire  _T_261; // @[Shift.scala 16:24]
  wire  _T_263; // @[Shift.scala 12:21]
  wire [2:0] _T_264; // @[Shift.scala 64:52]
  wire [10:0] _T_266; // @[Cat.scala 29:58]
  wire [10:0] _T_267; // @[Shift.scala 64:27]
  wire [2:0] _T_268; // @[Shift.scala 66:70]
  wire  _T_269; // @[Shift.scala 12:21]
  wire [6:0] _T_270; // @[Shift.scala 64:52]
  wire [10:0] _T_272; // @[Cat.scala 29:58]
  wire [10:0] _T_273; // @[Shift.scala 64:27]
  wire [1:0] _T_274; // @[Shift.scala 66:70]
  wire  _T_275; // @[Shift.scala 12:21]
  wire [8:0] _T_276; // @[Shift.scala 64:52]
  wire [10:0] _T_278; // @[Cat.scala 29:58]
  wire [10:0] _T_279; // @[Shift.scala 64:27]
  wire  _T_280; // @[Shift.scala 66:70]
  wire [9:0] _T_282; // @[Shift.scala 64:52]
  wire [10:0] _T_283; // @[Cat.scala 29:58]
  wire [10:0] _T_284; // @[Shift.scala 64:27]
  wire [10:0] _T_285; // @[Shift.scala 16:10]
  wire  _T_286; // @[convert.scala 23:34]
  wire [9:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_288; // @[convert.scala 25:26]
  wire [3:0] _T_290; // @[convert.scala 25:42]
  wire  _T_293; // @[convert.scala 26:67]
  wire  _T_294; // @[convert.scala 26:51]
  wire [5:0] _T_295; // @[Cat.scala 29:58]
  wire [12:0] _T_297; // @[convert.scala 29:56]
  wire  _T_298; // @[convert.scala 29:60]
  wire  _T_299; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_302; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [5:0] decB_scale; // @[convert.scala 32:24]
  wire  _T_311; // @[convert.scala 18:24]
  wire  _T_312; // @[convert.scala 18:40]
  wire  _T_313; // @[convert.scala 18:36]
  wire [11:0] _T_314; // @[convert.scala 19:24]
  wire [11:0] _T_315; // @[convert.scala 19:43]
  wire [11:0] _T_316; // @[convert.scala 19:39]
  wire [7:0] _T_317; // @[LZD.scala 43:32]
  wire [3:0] _T_318; // @[LZD.scala 43:32]
  wire [1:0] _T_319; // @[LZD.scala 43:32]
  wire  _T_320; // @[LZD.scala 39:14]
  wire  _T_321; // @[LZD.scala 39:21]
  wire  _T_322; // @[LZD.scala 39:30]
  wire  _T_323; // @[LZD.scala 39:27]
  wire  _T_324; // @[LZD.scala 39:25]
  wire [1:0] _T_325; // @[Cat.scala 29:58]
  wire [1:0] _T_326; // @[LZD.scala 44:32]
  wire  _T_327; // @[LZD.scala 39:14]
  wire  _T_328; // @[LZD.scala 39:21]
  wire  _T_329; // @[LZD.scala 39:30]
  wire  _T_330; // @[LZD.scala 39:27]
  wire  _T_331; // @[LZD.scala 39:25]
  wire [1:0] _T_332; // @[Cat.scala 29:58]
  wire  _T_333; // @[Shift.scala 12:21]
  wire  _T_334; // @[Shift.scala 12:21]
  wire  _T_335; // @[LZD.scala 49:16]
  wire  _T_336; // @[LZD.scala 49:27]
  wire  _T_337; // @[LZD.scala 49:25]
  wire  _T_338; // @[LZD.scala 49:47]
  wire  _T_339; // @[LZD.scala 49:59]
  wire  _T_340; // @[LZD.scala 49:35]
  wire [2:0] _T_342; // @[Cat.scala 29:58]
  wire [3:0] _T_343; // @[LZD.scala 44:32]
  wire [1:0] _T_344; // @[LZD.scala 43:32]
  wire  _T_345; // @[LZD.scala 39:14]
  wire  _T_346; // @[LZD.scala 39:21]
  wire  _T_347; // @[LZD.scala 39:30]
  wire  _T_348; // @[LZD.scala 39:27]
  wire  _T_349; // @[LZD.scala 39:25]
  wire [1:0] _T_350; // @[Cat.scala 29:58]
  wire [1:0] _T_351; // @[LZD.scala 44:32]
  wire  _T_352; // @[LZD.scala 39:14]
  wire  _T_353; // @[LZD.scala 39:21]
  wire  _T_354; // @[LZD.scala 39:30]
  wire  _T_355; // @[LZD.scala 39:27]
  wire  _T_356; // @[LZD.scala 39:25]
  wire [1:0] _T_357; // @[Cat.scala 29:58]
  wire  _T_358; // @[Shift.scala 12:21]
  wire  _T_359; // @[Shift.scala 12:21]
  wire  _T_360; // @[LZD.scala 49:16]
  wire  _T_361; // @[LZD.scala 49:27]
  wire  _T_362; // @[LZD.scala 49:25]
  wire  _T_363; // @[LZD.scala 49:47]
  wire  _T_364; // @[LZD.scala 49:59]
  wire  _T_365; // @[LZD.scala 49:35]
  wire [2:0] _T_367; // @[Cat.scala 29:58]
  wire  _T_368; // @[Shift.scala 12:21]
  wire  _T_369; // @[Shift.scala 12:21]
  wire  _T_370; // @[LZD.scala 49:16]
  wire  _T_371; // @[LZD.scala 49:27]
  wire  _T_372; // @[LZD.scala 49:25]
  wire [1:0] _T_373; // @[LZD.scala 49:47]
  wire [1:0] _T_374; // @[LZD.scala 49:59]
  wire [1:0] _T_375; // @[LZD.scala 49:35]
  wire [3:0] _T_377; // @[Cat.scala 29:58]
  wire [3:0] _T_378; // @[LZD.scala 44:32]
  wire [1:0] _T_379; // @[LZD.scala 43:32]
  wire  _T_380; // @[LZD.scala 39:14]
  wire  _T_381; // @[LZD.scala 39:21]
  wire  _T_382; // @[LZD.scala 39:30]
  wire  _T_383; // @[LZD.scala 39:27]
  wire  _T_384; // @[LZD.scala 39:25]
  wire [1:0] _T_385; // @[Cat.scala 29:58]
  wire [1:0] _T_386; // @[LZD.scala 44:32]
  wire  _T_387; // @[LZD.scala 39:14]
  wire  _T_388; // @[LZD.scala 39:21]
  wire  _T_389; // @[LZD.scala 39:30]
  wire  _T_390; // @[LZD.scala 39:27]
  wire  _T_391; // @[LZD.scala 39:25]
  wire [1:0] _T_392; // @[Cat.scala 29:58]
  wire  _T_393; // @[Shift.scala 12:21]
  wire  _T_394; // @[Shift.scala 12:21]
  wire  _T_395; // @[LZD.scala 49:16]
  wire  _T_396; // @[LZD.scala 49:27]
  wire  _T_397; // @[LZD.scala 49:25]
  wire  _T_398; // @[LZD.scala 49:47]
  wire  _T_399; // @[LZD.scala 49:59]
  wire  _T_400; // @[LZD.scala 49:35]
  wire [2:0] _T_402; // @[Cat.scala 29:58]
  wire  _T_403; // @[Shift.scala 12:21]
  wire [2:0] _T_405; // @[LZD.scala 55:32]
  wire [2:0] _T_406; // @[LZD.scala 55:20]
  wire [3:0] _T_407; // @[Cat.scala 29:58]
  wire [3:0] _T_408; // @[convert.scala 21:22]
  wire [10:0] _T_409; // @[convert.scala 22:36]
  wire  _T_410; // @[Shift.scala 16:24]
  wire  _T_412; // @[Shift.scala 12:21]
  wire [2:0] _T_413; // @[Shift.scala 64:52]
  wire [10:0] _T_415; // @[Cat.scala 29:58]
  wire [10:0] _T_416; // @[Shift.scala 64:27]
  wire [2:0] _T_417; // @[Shift.scala 66:70]
  wire  _T_418; // @[Shift.scala 12:21]
  wire [6:0] _T_419; // @[Shift.scala 64:52]
  wire [10:0] _T_421; // @[Cat.scala 29:58]
  wire [10:0] _T_422; // @[Shift.scala 64:27]
  wire [1:0] _T_423; // @[Shift.scala 66:70]
  wire  _T_424; // @[Shift.scala 12:21]
  wire [8:0] _T_425; // @[Shift.scala 64:52]
  wire [10:0] _T_427; // @[Cat.scala 29:58]
  wire [10:0] _T_428; // @[Shift.scala 64:27]
  wire  _T_429; // @[Shift.scala 66:70]
  wire [9:0] _T_431; // @[Shift.scala 64:52]
  wire [10:0] _T_432; // @[Cat.scala 29:58]
  wire [10:0] _T_433; // @[Shift.scala 64:27]
  wire [10:0] _T_434; // @[Shift.scala 16:10]
  wire  _T_435; // @[convert.scala 23:34]
  wire [9:0] decC_fraction; // @[convert.scala 24:34]
  wire  _T_437; // @[convert.scala 25:26]
  wire [3:0] _T_439; // @[convert.scala 25:42]
  wire  _T_442; // @[convert.scala 26:67]
  wire  _T_443; // @[convert.scala 26:51]
  wire [5:0] _T_444; // @[Cat.scala 29:58]
  wire [12:0] _T_446; // @[convert.scala 29:56]
  wire  _T_447; // @[convert.scala 29:60]
  wire  _T_448; // @[convert.scala 29:41]
  wire  decC_isNaR; // @[convert.scala 29:39]
  wire  _T_451; // @[convert.scala 30:19]
  wire  decC_isZero; // @[convert.scala 30:41]
  wire [5:0] decC_scale; // @[convert.scala 32:24]
  wire  _T_459; // @[PositFMA.scala 58:30]
  wire  outIsNaR; // @[PositFMA.scala 58:44]
  wire  _T_460; // @[PositFMA.scala 59:34]
  wire  _T_461; // @[PositFMA.scala 59:47]
  wire  _T_462; // @[PositFMA.scala 59:45]
  wire [11:0] _T_464; // @[Cat.scala 29:58]
  wire [11:0] sigA; // @[PositFMA.scala 59:76]
  wire  _T_465; // @[PositFMA.scala 60:34]
  wire  _T_466; // @[PositFMA.scala 60:47]
  wire  _T_467; // @[PositFMA.scala 60:45]
  wire [11:0] _T_469; // @[Cat.scala 29:58]
  wire [11:0] sigB; // @[PositFMA.scala 60:76]
  wire [23:0] _T_470; // @[PositFMA.scala 61:25]
  wire [23:0] sigP; // @[PositFMA.scala 61:33]
  wire [1:0] head2; // @[PositFMA.scala 62:28]
  wire  _T_471; // @[PositFMA.scala 63:31]
  wire  _T_472; // @[PositFMA.scala 63:25]
  wire  _T_473; // @[PositFMA.scala 63:42]
  wire  addTwo; // @[PositFMA.scala 63:35]
  wire  _T_474; // @[PositFMA.scala 65:23]
  wire  _T_475; // @[PositFMA.scala 65:49]
  wire  addOne; // @[PositFMA.scala 65:43]
  wire [1:0] _T_476; // @[Cat.scala 29:58]
  wire [2:0] expBias; // @[PositFMA.scala 66:39]
  wire  mulSign; // @[PositFMA.scala 67:28]
  wire [6:0] _T_477; // @[PositFMA.scala 69:30]
  wire [6:0] _GEN_12; // @[PositFMA.scala 69:44]
  wire [6:0] _T_479; // @[PositFMA.scala 69:44]
  wire [6:0] mulScale; // @[PositFMA.scala 69:44]
  wire [21:0] _T_480; // @[PositFMA.scala 72:29]
  wire [20:0] _T_481; // @[PositFMA.scala 73:29]
  wire [21:0] _T_482; // @[PositFMA.scala 73:48]
  wire [21:0] mulSigTmp; // @[PositFMA.scala 70:22]
  wire  _T_484; // @[PositFMA.scala 77:39]
  wire  _T_485; // @[PositFMA.scala 77:43]
  wire [20:0] _T_486; // @[PositFMA.scala 78:39]
  wire [22:0] mulSig; // @[Cat.scala 29:58]
  reg  outIsNaR_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg [22:0] mulSig_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg [9:0] addFrac_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [6:0] mulScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [5:0] addScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  addSign_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  addZero_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  inValid_phase2; // @[Valid.scala 117:22]
  reg [31:0] _RAND_7;
  wire  _T_512; // @[PositFMA.scala 107:29]
  wire  _T_513; // @[PositFMA.scala 107:47]
  wire  _T_514; // @[PositFMA.scala 107:45]
  wire [22:0] extAddSig; // @[Cat.scala 29:58]
  wire [6:0] _GEN_13; // @[PositFMA.scala 111:39]
  wire  mulGreater; // @[PositFMA.scala 111:39]
  wire [6:0] greaterScale; // @[PositFMA.scala 112:26]
  wire [6:0] smallerScale; // @[PositFMA.scala 113:26]
  wire [6:0] _T_518; // @[PositFMA.scala 114:36]
  wire [6:0] scaleDiff; // @[PositFMA.scala 114:36]
  wire [22:0] greaterSig; // @[PositFMA.scala 115:26]
  wire [22:0] smallerSigTmp; // @[PositFMA.scala 116:26]
  wire [6:0] _T_519; // @[PositFMA.scala 117:69]
  wire  _T_520; // @[Shift.scala 39:24]
  wire [4:0] _T_521; // @[Shift.scala 40:44]
  wire [6:0] _T_522; // @[Shift.scala 90:30]
  wire [15:0] _T_523; // @[Shift.scala 90:48]
  wire  _T_524; // @[Shift.scala 90:57]
  wire [6:0] _GEN_14; // @[Shift.scala 90:39]
  wire [6:0] _T_525; // @[Shift.scala 90:39]
  wire  _T_526; // @[Shift.scala 12:21]
  wire  _T_527; // @[Shift.scala 12:21]
  wire [15:0] _T_529; // @[Bitwise.scala 71:12]
  wire [22:0] _T_530; // @[Cat.scala 29:58]
  wire [22:0] _T_531; // @[Shift.scala 91:22]
  wire [3:0] _T_532; // @[Shift.scala 92:77]
  wire [14:0] _T_533; // @[Shift.scala 90:30]
  wire [7:0] _T_534; // @[Shift.scala 90:48]
  wire  _T_535; // @[Shift.scala 90:57]
  wire [14:0] _GEN_15; // @[Shift.scala 90:39]
  wire [14:0] _T_536; // @[Shift.scala 90:39]
  wire  _T_537; // @[Shift.scala 12:21]
  wire  _T_538; // @[Shift.scala 12:21]
  wire [7:0] _T_540; // @[Bitwise.scala 71:12]
  wire [22:0] _T_541; // @[Cat.scala 29:58]
  wire [22:0] _T_542; // @[Shift.scala 91:22]
  wire [2:0] _T_543; // @[Shift.scala 92:77]
  wire [18:0] _T_544; // @[Shift.scala 90:30]
  wire [3:0] _T_545; // @[Shift.scala 90:48]
  wire  _T_546; // @[Shift.scala 90:57]
  wire [18:0] _GEN_16; // @[Shift.scala 90:39]
  wire [18:0] _T_547; // @[Shift.scala 90:39]
  wire  _T_548; // @[Shift.scala 12:21]
  wire  _T_549; // @[Shift.scala 12:21]
  wire [3:0] _T_551; // @[Bitwise.scala 71:12]
  wire [22:0] _T_552; // @[Cat.scala 29:58]
  wire [22:0] _T_553; // @[Shift.scala 91:22]
  wire [1:0] _T_554; // @[Shift.scala 92:77]
  wire [20:0] _T_555; // @[Shift.scala 90:30]
  wire [1:0] _T_556; // @[Shift.scala 90:48]
  wire  _T_557; // @[Shift.scala 90:57]
  wire [20:0] _GEN_17; // @[Shift.scala 90:39]
  wire [20:0] _T_558; // @[Shift.scala 90:39]
  wire  _T_559; // @[Shift.scala 12:21]
  wire  _T_560; // @[Shift.scala 12:21]
  wire [1:0] _T_562; // @[Bitwise.scala 71:12]
  wire [22:0] _T_563; // @[Cat.scala 29:58]
  wire [22:0] _T_564; // @[Shift.scala 91:22]
  wire  _T_565; // @[Shift.scala 92:77]
  wire [21:0] _T_566; // @[Shift.scala 90:30]
  wire  _T_567; // @[Shift.scala 90:48]
  wire [21:0] _GEN_18; // @[Shift.scala 90:39]
  wire [21:0] _T_569; // @[Shift.scala 90:39]
  wire  _T_571; // @[Shift.scala 12:21]
  wire [22:0] _T_572; // @[Cat.scala 29:58]
  wire [22:0] _T_573; // @[Shift.scala 91:22]
  wire [22:0] _T_576; // @[Bitwise.scala 71:12]
  wire [22:0] smallerSig; // @[Shift.scala 39:10]
  wire [23:0] rawSumSig; // @[PositFMA.scala 118:34]
  wire  _T_577; // @[PositFMA.scala 119:42]
  wire  _T_578; // @[PositFMA.scala 119:46]
  wire  _T_579; // @[PositFMA.scala 119:79]
  wire  sumSign; // @[PositFMA.scala 119:63]
  wire [22:0] _T_581; // @[PositFMA.scala 120:50]
  wire [23:0] signSumSig; // @[Cat.scala 29:58]
  wire [22:0] _T_582; // @[PositFMA.scala 124:33]
  wire [22:0] _T_583; // @[PositFMA.scala 124:68]
  wire [22:0] sumXor; // @[PositFMA.scala 124:51]
  wire [15:0] _T_584; // @[LZD.scala 43:32]
  wire [7:0] _T_585; // @[LZD.scala 43:32]
  wire [3:0] _T_586; // @[LZD.scala 43:32]
  wire [1:0] _T_587; // @[LZD.scala 43:32]
  wire  _T_588; // @[LZD.scala 39:14]
  wire  _T_589; // @[LZD.scala 39:21]
  wire  _T_590; // @[LZD.scala 39:30]
  wire  _T_591; // @[LZD.scala 39:27]
  wire  _T_592; // @[LZD.scala 39:25]
  wire [1:0] _T_593; // @[Cat.scala 29:58]
  wire [1:0] _T_594; // @[LZD.scala 44:32]
  wire  _T_595; // @[LZD.scala 39:14]
  wire  _T_596; // @[LZD.scala 39:21]
  wire  _T_597; // @[LZD.scala 39:30]
  wire  _T_598; // @[LZD.scala 39:27]
  wire  _T_599; // @[LZD.scala 39:25]
  wire [1:0] _T_600; // @[Cat.scala 29:58]
  wire  _T_601; // @[Shift.scala 12:21]
  wire  _T_602; // @[Shift.scala 12:21]
  wire  _T_603; // @[LZD.scala 49:16]
  wire  _T_604; // @[LZD.scala 49:27]
  wire  _T_605; // @[LZD.scala 49:25]
  wire  _T_606; // @[LZD.scala 49:47]
  wire  _T_607; // @[LZD.scala 49:59]
  wire  _T_608; // @[LZD.scala 49:35]
  wire [2:0] _T_610; // @[Cat.scala 29:58]
  wire [3:0] _T_611; // @[LZD.scala 44:32]
  wire [1:0] _T_612; // @[LZD.scala 43:32]
  wire  _T_613; // @[LZD.scala 39:14]
  wire  _T_614; // @[LZD.scala 39:21]
  wire  _T_615; // @[LZD.scala 39:30]
  wire  _T_616; // @[LZD.scala 39:27]
  wire  _T_617; // @[LZD.scala 39:25]
  wire [1:0] _T_618; // @[Cat.scala 29:58]
  wire [1:0] _T_619; // @[LZD.scala 44:32]
  wire  _T_620; // @[LZD.scala 39:14]
  wire  _T_621; // @[LZD.scala 39:21]
  wire  _T_622; // @[LZD.scala 39:30]
  wire  _T_623; // @[LZD.scala 39:27]
  wire  _T_624; // @[LZD.scala 39:25]
  wire [1:0] _T_625; // @[Cat.scala 29:58]
  wire  _T_626; // @[Shift.scala 12:21]
  wire  _T_627; // @[Shift.scala 12:21]
  wire  _T_628; // @[LZD.scala 49:16]
  wire  _T_629; // @[LZD.scala 49:27]
  wire  _T_630; // @[LZD.scala 49:25]
  wire  _T_631; // @[LZD.scala 49:47]
  wire  _T_632; // @[LZD.scala 49:59]
  wire  _T_633; // @[LZD.scala 49:35]
  wire [2:0] _T_635; // @[Cat.scala 29:58]
  wire  _T_636; // @[Shift.scala 12:21]
  wire  _T_637; // @[Shift.scala 12:21]
  wire  _T_638; // @[LZD.scala 49:16]
  wire  _T_639; // @[LZD.scala 49:27]
  wire  _T_640; // @[LZD.scala 49:25]
  wire [1:0] _T_641; // @[LZD.scala 49:47]
  wire [1:0] _T_642; // @[LZD.scala 49:59]
  wire [1:0] _T_643; // @[LZD.scala 49:35]
  wire [3:0] _T_645; // @[Cat.scala 29:58]
  wire [7:0] _T_646; // @[LZD.scala 44:32]
  wire [3:0] _T_647; // @[LZD.scala 43:32]
  wire [1:0] _T_648; // @[LZD.scala 43:32]
  wire  _T_649; // @[LZD.scala 39:14]
  wire  _T_650; // @[LZD.scala 39:21]
  wire  _T_651; // @[LZD.scala 39:30]
  wire  _T_652; // @[LZD.scala 39:27]
  wire  _T_653; // @[LZD.scala 39:25]
  wire [1:0] _T_654; // @[Cat.scala 29:58]
  wire [1:0] _T_655; // @[LZD.scala 44:32]
  wire  _T_656; // @[LZD.scala 39:14]
  wire  _T_657; // @[LZD.scala 39:21]
  wire  _T_658; // @[LZD.scala 39:30]
  wire  _T_659; // @[LZD.scala 39:27]
  wire  _T_660; // @[LZD.scala 39:25]
  wire [1:0] _T_661; // @[Cat.scala 29:58]
  wire  _T_662; // @[Shift.scala 12:21]
  wire  _T_663; // @[Shift.scala 12:21]
  wire  _T_664; // @[LZD.scala 49:16]
  wire  _T_665; // @[LZD.scala 49:27]
  wire  _T_666; // @[LZD.scala 49:25]
  wire  _T_667; // @[LZD.scala 49:47]
  wire  _T_668; // @[LZD.scala 49:59]
  wire  _T_669; // @[LZD.scala 49:35]
  wire [2:0] _T_671; // @[Cat.scala 29:58]
  wire [3:0] _T_672; // @[LZD.scala 44:32]
  wire [1:0] _T_673; // @[LZD.scala 43:32]
  wire  _T_674; // @[LZD.scala 39:14]
  wire  _T_675; // @[LZD.scala 39:21]
  wire  _T_676; // @[LZD.scala 39:30]
  wire  _T_677; // @[LZD.scala 39:27]
  wire  _T_678; // @[LZD.scala 39:25]
  wire [1:0] _T_679; // @[Cat.scala 29:58]
  wire [1:0] _T_680; // @[LZD.scala 44:32]
  wire  _T_681; // @[LZD.scala 39:14]
  wire  _T_682; // @[LZD.scala 39:21]
  wire  _T_683; // @[LZD.scala 39:30]
  wire  _T_684; // @[LZD.scala 39:27]
  wire  _T_685; // @[LZD.scala 39:25]
  wire [1:0] _T_686; // @[Cat.scala 29:58]
  wire  _T_687; // @[Shift.scala 12:21]
  wire  _T_688; // @[Shift.scala 12:21]
  wire  _T_689; // @[LZD.scala 49:16]
  wire  _T_690; // @[LZD.scala 49:27]
  wire  _T_691; // @[LZD.scala 49:25]
  wire  _T_692; // @[LZD.scala 49:47]
  wire  _T_693; // @[LZD.scala 49:59]
  wire  _T_694; // @[LZD.scala 49:35]
  wire [2:0] _T_696; // @[Cat.scala 29:58]
  wire  _T_697; // @[Shift.scala 12:21]
  wire  _T_698; // @[Shift.scala 12:21]
  wire  _T_699; // @[LZD.scala 49:16]
  wire  _T_700; // @[LZD.scala 49:27]
  wire  _T_701; // @[LZD.scala 49:25]
  wire [1:0] _T_702; // @[LZD.scala 49:47]
  wire [1:0] _T_703; // @[LZD.scala 49:59]
  wire [1:0] _T_704; // @[LZD.scala 49:35]
  wire [3:0] _T_706; // @[Cat.scala 29:58]
  wire  _T_707; // @[Shift.scala 12:21]
  wire  _T_708; // @[Shift.scala 12:21]
  wire  _T_709; // @[LZD.scala 49:16]
  wire  _T_710; // @[LZD.scala 49:27]
  wire  _T_711; // @[LZD.scala 49:25]
  wire [2:0] _T_712; // @[LZD.scala 49:47]
  wire [2:0] _T_713; // @[LZD.scala 49:59]
  wire [2:0] _T_714; // @[LZD.scala 49:35]
  wire [4:0] _T_716; // @[Cat.scala 29:58]
  wire [6:0] _T_717; // @[LZD.scala 44:32]
  wire [3:0] _T_718; // @[LZD.scala 43:32]
  wire [1:0] _T_719; // @[LZD.scala 43:32]
  wire  _T_720; // @[LZD.scala 39:14]
  wire  _T_721; // @[LZD.scala 39:21]
  wire  _T_722; // @[LZD.scala 39:30]
  wire  _T_723; // @[LZD.scala 39:27]
  wire  _T_724; // @[LZD.scala 39:25]
  wire [1:0] _T_725; // @[Cat.scala 29:58]
  wire [1:0] _T_726; // @[LZD.scala 44:32]
  wire  _T_727; // @[LZD.scala 39:14]
  wire  _T_728; // @[LZD.scala 39:21]
  wire  _T_729; // @[LZD.scala 39:30]
  wire  _T_730; // @[LZD.scala 39:27]
  wire  _T_731; // @[LZD.scala 39:25]
  wire [1:0] _T_732; // @[Cat.scala 29:58]
  wire  _T_733; // @[Shift.scala 12:21]
  wire  _T_734; // @[Shift.scala 12:21]
  wire  _T_735; // @[LZD.scala 49:16]
  wire  _T_736; // @[LZD.scala 49:27]
  wire  _T_737; // @[LZD.scala 49:25]
  wire  _T_738; // @[LZD.scala 49:47]
  wire  _T_739; // @[LZD.scala 49:59]
  wire  _T_740; // @[LZD.scala 49:35]
  wire [2:0] _T_742; // @[Cat.scala 29:58]
  wire [2:0] _T_743; // @[LZD.scala 44:32]
  wire [1:0] _T_744; // @[LZD.scala 43:32]
  wire  _T_745; // @[LZD.scala 39:14]
  wire  _T_746; // @[LZD.scala 39:21]
  wire  _T_747; // @[LZD.scala 39:30]
  wire  _T_748; // @[LZD.scala 39:27]
  wire  _T_749; // @[LZD.scala 39:25]
  wire [1:0] _T_750; // @[Cat.scala 29:58]
  wire  _T_751; // @[LZD.scala 44:32]
  wire  _T_753; // @[Shift.scala 12:21]
  wire  _T_755; // @[LZD.scala 55:32]
  wire  _T_756; // @[LZD.scala 55:20]
  wire [1:0] _T_757; // @[Cat.scala 29:58]
  wire  _T_758; // @[Shift.scala 12:21]
  wire [1:0] _T_760; // @[LZD.scala 55:32]
  wire [1:0] _T_761; // @[LZD.scala 55:20]
  wire  _T_763; // @[Shift.scala 12:21]
  wire [3:0] _T_765; // @[Cat.scala 29:58]
  wire [3:0] _T_766; // @[LZD.scala 55:32]
  wire [3:0] _T_767; // @[LZD.scala 55:20]
  wire [4:0] sumLZD; // @[Cat.scala 29:58]
  wire [4:0] shiftValue; // @[PositFMA.scala 126:24]
  wire [21:0] _T_768; // @[PositFMA.scala 127:38]
  wire  _T_769; // @[Shift.scala 16:24]
  wire  _T_771; // @[Shift.scala 12:21]
  wire [5:0] _T_772; // @[Shift.scala 64:52]
  wire [21:0] _T_774; // @[Cat.scala 29:58]
  wire [21:0] _T_775; // @[Shift.scala 64:27]
  wire [3:0] _T_776; // @[Shift.scala 66:70]
  wire  _T_777; // @[Shift.scala 12:21]
  wire [13:0] _T_778; // @[Shift.scala 64:52]
  wire [21:0] _T_780; // @[Cat.scala 29:58]
  wire [21:0] _T_781; // @[Shift.scala 64:27]
  wire [2:0] _T_782; // @[Shift.scala 66:70]
  wire  _T_783; // @[Shift.scala 12:21]
  wire [17:0] _T_784; // @[Shift.scala 64:52]
  wire [21:0] _T_786; // @[Cat.scala 29:58]
  wire [21:0] _T_787; // @[Shift.scala 64:27]
  wire [1:0] _T_788; // @[Shift.scala 66:70]
  wire  _T_789; // @[Shift.scala 12:21]
  wire [19:0] _T_790; // @[Shift.scala 64:52]
  wire [21:0] _T_792; // @[Cat.scala 29:58]
  wire [21:0] _T_793; // @[Shift.scala 64:27]
  wire  _T_794; // @[Shift.scala 66:70]
  wire [20:0] _T_796; // @[Shift.scala 64:52]
  wire [21:0] _T_797; // @[Cat.scala 29:58]
  wire [21:0] _T_798; // @[Shift.scala 64:27]
  wire [21:0] normalFracTmp; // @[Shift.scala 16:10]
  wire [6:0] _T_800; // @[PositFMA.scala 130:36]
  wire [6:0] _T_801; // @[PositFMA.scala 130:36]
  wire [5:0] _T_802; // @[Cat.scala 29:58]
  wire [5:0] _T_803; // @[PositFMA.scala 130:61]
  wire [6:0] _GEN_19; // @[PositFMA.scala 130:42]
  wire [6:0] _T_805; // @[PositFMA.scala 130:42]
  wire [6:0] sumScale; // @[PositFMA.scala 130:42]
  wire [9:0] sumFrac; // @[PositFMA.scala 131:41]
  wire [11:0] grsTmp; // @[PositFMA.scala 134:41]
  wire [1:0] _T_806; // @[PositFMA.scala 137:40]
  wire [9:0] _T_807; // @[PositFMA.scala 137:56]
  wire  _T_808; // @[PositFMA.scala 137:60]
  wire  underflow; // @[PositFMA.scala 144:32]
  wire  overflow; // @[PositFMA.scala 145:32]
  wire  _T_809; // @[PositFMA.scala 154:32]
  wire  decF_isZero; // @[PositFMA.scala 154:20]
  wire [6:0] _T_811; // @[Mux.scala 87:16]
  wire [6:0] _T_812; // @[Mux.scala 87:16]
  wire [5:0] _GEN_20; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  wire [5:0] decF_scale; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  wire  _T_813; // @[convert.scala 46:61]
  wire  _T_814; // @[convert.scala 46:52]
  wire  _T_816; // @[convert.scala 46:42]
  wire [4:0] _T_817; // @[convert.scala 48:34]
  wire  _T_818; // @[convert.scala 49:36]
  wire [4:0] _T_820; // @[convert.scala 50:36]
  wire [4:0] _T_821; // @[convert.scala 50:36]
  wire [4:0] _T_822; // @[convert.scala 50:28]
  wire  _T_823; // @[convert.scala 51:31]
  wire  _T_824; // @[convert.scala 52:43]
  wire [15:0] _T_828; // @[Cat.scala 29:58]
  wire [4:0] _T_829; // @[Shift.scala 39:17]
  wire  _T_830; // @[Shift.scala 39:24]
  wire [3:0] _T_831; // @[Shift.scala 40:44]
  wire [7:0] _T_832; // @[Shift.scala 90:30]
  wire [7:0] _T_833; // @[Shift.scala 90:48]
  wire  _T_834; // @[Shift.scala 90:57]
  wire [7:0] _GEN_21; // @[Shift.scala 90:39]
  wire [7:0] _T_835; // @[Shift.scala 90:39]
  wire  _T_836; // @[Shift.scala 12:21]
  wire  _T_837; // @[Shift.scala 12:21]
  wire [7:0] _T_839; // @[Bitwise.scala 71:12]
  wire [15:0] _T_840; // @[Cat.scala 29:58]
  wire [15:0] _T_841; // @[Shift.scala 91:22]
  wire [2:0] _T_842; // @[Shift.scala 92:77]
  wire [11:0] _T_843; // @[Shift.scala 90:30]
  wire [3:0] _T_844; // @[Shift.scala 90:48]
  wire  _T_845; // @[Shift.scala 90:57]
  wire [11:0] _GEN_22; // @[Shift.scala 90:39]
  wire [11:0] _T_846; // @[Shift.scala 90:39]
  wire  _T_847; // @[Shift.scala 12:21]
  wire  _T_848; // @[Shift.scala 12:21]
  wire [3:0] _T_850; // @[Bitwise.scala 71:12]
  wire [15:0] _T_851; // @[Cat.scala 29:58]
  wire [15:0] _T_852; // @[Shift.scala 91:22]
  wire [1:0] _T_853; // @[Shift.scala 92:77]
  wire [13:0] _T_854; // @[Shift.scala 90:30]
  wire [1:0] _T_855; // @[Shift.scala 90:48]
  wire  _T_856; // @[Shift.scala 90:57]
  wire [13:0] _GEN_23; // @[Shift.scala 90:39]
  wire [13:0] _T_857; // @[Shift.scala 90:39]
  wire  _T_858; // @[Shift.scala 12:21]
  wire  _T_859; // @[Shift.scala 12:21]
  wire [1:0] _T_861; // @[Bitwise.scala 71:12]
  wire [15:0] _T_862; // @[Cat.scala 29:58]
  wire [15:0] _T_863; // @[Shift.scala 91:22]
  wire  _T_864; // @[Shift.scala 92:77]
  wire [14:0] _T_865; // @[Shift.scala 90:30]
  wire  _T_866; // @[Shift.scala 90:48]
  wire [14:0] _GEN_24; // @[Shift.scala 90:39]
  wire [14:0] _T_868; // @[Shift.scala 90:39]
  wire  _T_870; // @[Shift.scala 12:21]
  wire [15:0] _T_871; // @[Cat.scala 29:58]
  wire [15:0] _T_872; // @[Shift.scala 91:22]
  wire [15:0] _T_875; // @[Bitwise.scala 71:12]
  wire [15:0] _T_876; // @[Shift.scala 39:10]
  wire  _T_877; // @[convert.scala 55:31]
  wire  _T_878; // @[convert.scala 56:31]
  wire  _T_879; // @[convert.scala 57:31]
  wire  _T_880; // @[convert.scala 58:31]
  wire [12:0] _T_881; // @[convert.scala 59:69]
  wire  _T_882; // @[convert.scala 59:81]
  wire  _T_883; // @[convert.scala 59:50]
  wire  _T_885; // @[convert.scala 60:81]
  wire  _T_886; // @[convert.scala 61:44]
  wire  _T_887; // @[convert.scala 61:52]
  wire  _T_888; // @[convert.scala 61:36]
  wire  _T_889; // @[convert.scala 62:63]
  wire  _T_890; // @[convert.scala 62:103]
  wire  _T_891; // @[convert.scala 62:60]
  wire [12:0] _GEN_25; // @[convert.scala 63:56]
  wire [12:0] _T_894; // @[convert.scala 63:56]
  wire [13:0] _T_895; // @[Cat.scala 29:58]
  reg  _T_899; // @[Valid.scala 117:22]
  reg [31:0] _RAND_8;
  reg [13:0] _T_903; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  assign _T = io_fmaOp[1]; // @[PositFMA.scala 47:36]
  assign _T_2 = _T ? 14'h3fff : 14'h0; // @[Bitwise.scala 71:12]
  assign _T_3 = _T_2 ^ io_A; // @[PositFMA.scala 47:41]
  assign _GEN_10 = {{13'd0}, _T}; // @[PositFMA.scala 47:49]
  assign realA = _T_3 + _GEN_10; // @[PositFMA.scala 47:49]
  assign _T_6 = io_fmaOp[0]; // @[PositFMA.scala 48:36]
  assign _T_8 = _T_6 ? 14'h3fff : 14'h0; // @[Bitwise.scala 71:12]
  assign _T_9 = _T_8 ^ io_C; // @[PositFMA.scala 48:41]
  assign _GEN_11 = {{13'd0}, _T_6}; // @[PositFMA.scala 48:49]
  assign realC = _T_9 + _GEN_11; // @[PositFMA.scala 48:49]
  assign _T_13 = realA[13]; // @[convert.scala 18:24]
  assign _T_14 = realA[12]; // @[convert.scala 18:40]
  assign _T_15 = _T_13 ^ _T_14; // @[convert.scala 18:36]
  assign _T_16 = realA[12:1]; // @[convert.scala 19:24]
  assign _T_17 = realA[11:0]; // @[convert.scala 19:43]
  assign _T_18 = _T_16 ^ _T_17; // @[convert.scala 19:39]
  assign _T_19 = _T_18[11:4]; // @[LZD.scala 43:32]
  assign _T_20 = _T_19[7:4]; // @[LZD.scala 43:32]
  assign _T_21 = _T_20[3:2]; // @[LZD.scala 43:32]
  assign _T_22 = _T_21 != 2'h0; // @[LZD.scala 39:14]
  assign _T_23 = _T_21[1]; // @[LZD.scala 39:21]
  assign _T_24 = _T_21[0]; // @[LZD.scala 39:30]
  assign _T_25 = ~ _T_24; // @[LZD.scala 39:27]
  assign _T_26 = _T_23 | _T_25; // @[LZD.scala 39:25]
  assign _T_27 = {_T_22,_T_26}; // @[Cat.scala 29:58]
  assign _T_28 = _T_20[1:0]; // @[LZD.scala 44:32]
  assign _T_29 = _T_28 != 2'h0; // @[LZD.scala 39:14]
  assign _T_30 = _T_28[1]; // @[LZD.scala 39:21]
  assign _T_31 = _T_28[0]; // @[LZD.scala 39:30]
  assign _T_32 = ~ _T_31; // @[LZD.scala 39:27]
  assign _T_33 = _T_30 | _T_32; // @[LZD.scala 39:25]
  assign _T_34 = {_T_29,_T_33}; // @[Cat.scala 29:58]
  assign _T_35 = _T_27[1]; // @[Shift.scala 12:21]
  assign _T_36 = _T_34[1]; // @[Shift.scala 12:21]
  assign _T_37 = _T_35 | _T_36; // @[LZD.scala 49:16]
  assign _T_38 = ~ _T_36; // @[LZD.scala 49:27]
  assign _T_39 = _T_35 | _T_38; // @[LZD.scala 49:25]
  assign _T_40 = _T_27[0:0]; // @[LZD.scala 49:47]
  assign _T_41 = _T_34[0:0]; // @[LZD.scala 49:59]
  assign _T_42 = _T_35 ? _T_40 : _T_41; // @[LZD.scala 49:35]
  assign _T_44 = {_T_37,_T_39,_T_42}; // @[Cat.scala 29:58]
  assign _T_45 = _T_19[3:0]; // @[LZD.scala 44:32]
  assign _T_46 = _T_45[3:2]; // @[LZD.scala 43:32]
  assign _T_47 = _T_46 != 2'h0; // @[LZD.scala 39:14]
  assign _T_48 = _T_46[1]; // @[LZD.scala 39:21]
  assign _T_49 = _T_46[0]; // @[LZD.scala 39:30]
  assign _T_50 = ~ _T_49; // @[LZD.scala 39:27]
  assign _T_51 = _T_48 | _T_50; // @[LZD.scala 39:25]
  assign _T_52 = {_T_47,_T_51}; // @[Cat.scala 29:58]
  assign _T_53 = _T_45[1:0]; // @[LZD.scala 44:32]
  assign _T_54 = _T_53 != 2'h0; // @[LZD.scala 39:14]
  assign _T_55 = _T_53[1]; // @[LZD.scala 39:21]
  assign _T_56 = _T_53[0]; // @[LZD.scala 39:30]
  assign _T_57 = ~ _T_56; // @[LZD.scala 39:27]
  assign _T_58 = _T_55 | _T_57; // @[LZD.scala 39:25]
  assign _T_59 = {_T_54,_T_58}; // @[Cat.scala 29:58]
  assign _T_60 = _T_52[1]; // @[Shift.scala 12:21]
  assign _T_61 = _T_59[1]; // @[Shift.scala 12:21]
  assign _T_62 = _T_60 | _T_61; // @[LZD.scala 49:16]
  assign _T_63 = ~ _T_61; // @[LZD.scala 49:27]
  assign _T_64 = _T_60 | _T_63; // @[LZD.scala 49:25]
  assign _T_65 = _T_52[0:0]; // @[LZD.scala 49:47]
  assign _T_66 = _T_59[0:0]; // @[LZD.scala 49:59]
  assign _T_67 = _T_60 ? _T_65 : _T_66; // @[LZD.scala 49:35]
  assign _T_69 = {_T_62,_T_64,_T_67}; // @[Cat.scala 29:58]
  assign _T_70 = _T_44[2]; // @[Shift.scala 12:21]
  assign _T_71 = _T_69[2]; // @[Shift.scala 12:21]
  assign _T_72 = _T_70 | _T_71; // @[LZD.scala 49:16]
  assign _T_73 = ~ _T_71; // @[LZD.scala 49:27]
  assign _T_74 = _T_70 | _T_73; // @[LZD.scala 49:25]
  assign _T_75 = _T_44[1:0]; // @[LZD.scala 49:47]
  assign _T_76 = _T_69[1:0]; // @[LZD.scala 49:59]
  assign _T_77 = _T_70 ? _T_75 : _T_76; // @[LZD.scala 49:35]
  assign _T_79 = {_T_72,_T_74,_T_77}; // @[Cat.scala 29:58]
  assign _T_80 = _T_18[3:0]; // @[LZD.scala 44:32]
  assign _T_81 = _T_80[3:2]; // @[LZD.scala 43:32]
  assign _T_82 = _T_81 != 2'h0; // @[LZD.scala 39:14]
  assign _T_83 = _T_81[1]; // @[LZD.scala 39:21]
  assign _T_84 = _T_81[0]; // @[LZD.scala 39:30]
  assign _T_85 = ~ _T_84; // @[LZD.scala 39:27]
  assign _T_86 = _T_83 | _T_85; // @[LZD.scala 39:25]
  assign _T_87 = {_T_82,_T_86}; // @[Cat.scala 29:58]
  assign _T_88 = _T_80[1:0]; // @[LZD.scala 44:32]
  assign _T_89 = _T_88 != 2'h0; // @[LZD.scala 39:14]
  assign _T_90 = _T_88[1]; // @[LZD.scala 39:21]
  assign _T_91 = _T_88[0]; // @[LZD.scala 39:30]
  assign _T_92 = ~ _T_91; // @[LZD.scala 39:27]
  assign _T_93 = _T_90 | _T_92; // @[LZD.scala 39:25]
  assign _T_94 = {_T_89,_T_93}; // @[Cat.scala 29:58]
  assign _T_95 = _T_87[1]; // @[Shift.scala 12:21]
  assign _T_96 = _T_94[1]; // @[Shift.scala 12:21]
  assign _T_97 = _T_95 | _T_96; // @[LZD.scala 49:16]
  assign _T_98 = ~ _T_96; // @[LZD.scala 49:27]
  assign _T_99 = _T_95 | _T_98; // @[LZD.scala 49:25]
  assign _T_100 = _T_87[0:0]; // @[LZD.scala 49:47]
  assign _T_101 = _T_94[0:0]; // @[LZD.scala 49:59]
  assign _T_102 = _T_95 ? _T_100 : _T_101; // @[LZD.scala 49:35]
  assign _T_104 = {_T_97,_T_99,_T_102}; // @[Cat.scala 29:58]
  assign _T_105 = _T_79[3]; // @[Shift.scala 12:21]
  assign _T_107 = _T_79[2:0]; // @[LZD.scala 55:32]
  assign _T_108 = _T_105 ? _T_107 : _T_104; // @[LZD.scala 55:20]
  assign _T_109 = {_T_105,_T_108}; // @[Cat.scala 29:58]
  assign _T_110 = ~ _T_109; // @[convert.scala 21:22]
  assign _T_111 = realA[10:0]; // @[convert.scala 22:36]
  assign _T_112 = _T_110 < 4'hb; // @[Shift.scala 16:24]
  assign _T_114 = _T_110[3]; // @[Shift.scala 12:21]
  assign _T_115 = _T_111[2:0]; // @[Shift.scala 64:52]
  assign _T_117 = {_T_115,8'h0}; // @[Cat.scala 29:58]
  assign _T_118 = _T_114 ? _T_117 : _T_111; // @[Shift.scala 64:27]
  assign _T_119 = _T_110[2:0]; // @[Shift.scala 66:70]
  assign _T_120 = _T_119[2]; // @[Shift.scala 12:21]
  assign _T_121 = _T_118[6:0]; // @[Shift.scala 64:52]
  assign _T_123 = {_T_121,4'h0}; // @[Cat.scala 29:58]
  assign _T_124 = _T_120 ? _T_123 : _T_118; // @[Shift.scala 64:27]
  assign _T_125 = _T_119[1:0]; // @[Shift.scala 66:70]
  assign _T_126 = _T_125[1]; // @[Shift.scala 12:21]
  assign _T_127 = _T_124[8:0]; // @[Shift.scala 64:52]
  assign _T_129 = {_T_127,2'h0}; // @[Cat.scala 29:58]
  assign _T_130 = _T_126 ? _T_129 : _T_124; // @[Shift.scala 64:27]
  assign _T_131 = _T_125[0:0]; // @[Shift.scala 66:70]
  assign _T_133 = _T_130[9:0]; // @[Shift.scala 64:52]
  assign _T_134 = {_T_133,1'h0}; // @[Cat.scala 29:58]
  assign _T_135 = _T_131 ? _T_134 : _T_130; // @[Shift.scala 64:27]
  assign _T_136 = _T_112 ? _T_135 : 11'h0; // @[Shift.scala 16:10]
  assign _T_137 = _T_136[10:10]; // @[convert.scala 23:34]
  assign decA_fraction = _T_136[9:0]; // @[convert.scala 24:34]
  assign _T_139 = _T_15 == 1'h0; // @[convert.scala 25:26]
  assign _T_141 = _T_15 ? _T_110 : _T_109; // @[convert.scala 25:42]
  assign _T_144 = ~ _T_137; // @[convert.scala 26:67]
  assign _T_145 = _T_13 ? _T_144 : _T_137; // @[convert.scala 26:51]
  assign _T_146 = {_T_139,_T_141,_T_145}; // @[Cat.scala 29:58]
  assign _T_148 = realA[12:0]; // @[convert.scala 29:56]
  assign _T_149 = _T_148 != 13'h0; // @[convert.scala 29:60]
  assign _T_150 = ~ _T_149; // @[convert.scala 29:41]
  assign decA_isNaR = _T_13 & _T_150; // @[convert.scala 29:39]
  assign _T_153 = _T_13 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_153 & _T_150; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_146); // @[convert.scala 32:24]
  assign _T_162 = io_B[13]; // @[convert.scala 18:24]
  assign _T_163 = io_B[12]; // @[convert.scala 18:40]
  assign _T_164 = _T_162 ^ _T_163; // @[convert.scala 18:36]
  assign _T_165 = io_B[12:1]; // @[convert.scala 19:24]
  assign _T_166 = io_B[11:0]; // @[convert.scala 19:43]
  assign _T_167 = _T_165 ^ _T_166; // @[convert.scala 19:39]
  assign _T_168 = _T_167[11:4]; // @[LZD.scala 43:32]
  assign _T_169 = _T_168[7:4]; // @[LZD.scala 43:32]
  assign _T_170 = _T_169[3:2]; // @[LZD.scala 43:32]
  assign _T_171 = _T_170 != 2'h0; // @[LZD.scala 39:14]
  assign _T_172 = _T_170[1]; // @[LZD.scala 39:21]
  assign _T_173 = _T_170[0]; // @[LZD.scala 39:30]
  assign _T_174 = ~ _T_173; // @[LZD.scala 39:27]
  assign _T_175 = _T_172 | _T_174; // @[LZD.scala 39:25]
  assign _T_176 = {_T_171,_T_175}; // @[Cat.scala 29:58]
  assign _T_177 = _T_169[1:0]; // @[LZD.scala 44:32]
  assign _T_178 = _T_177 != 2'h0; // @[LZD.scala 39:14]
  assign _T_179 = _T_177[1]; // @[LZD.scala 39:21]
  assign _T_180 = _T_177[0]; // @[LZD.scala 39:30]
  assign _T_181 = ~ _T_180; // @[LZD.scala 39:27]
  assign _T_182 = _T_179 | _T_181; // @[LZD.scala 39:25]
  assign _T_183 = {_T_178,_T_182}; // @[Cat.scala 29:58]
  assign _T_184 = _T_176[1]; // @[Shift.scala 12:21]
  assign _T_185 = _T_183[1]; // @[Shift.scala 12:21]
  assign _T_186 = _T_184 | _T_185; // @[LZD.scala 49:16]
  assign _T_187 = ~ _T_185; // @[LZD.scala 49:27]
  assign _T_188 = _T_184 | _T_187; // @[LZD.scala 49:25]
  assign _T_189 = _T_176[0:0]; // @[LZD.scala 49:47]
  assign _T_190 = _T_183[0:0]; // @[LZD.scala 49:59]
  assign _T_191 = _T_184 ? _T_189 : _T_190; // @[LZD.scala 49:35]
  assign _T_193 = {_T_186,_T_188,_T_191}; // @[Cat.scala 29:58]
  assign _T_194 = _T_168[3:0]; // @[LZD.scala 44:32]
  assign _T_195 = _T_194[3:2]; // @[LZD.scala 43:32]
  assign _T_196 = _T_195 != 2'h0; // @[LZD.scala 39:14]
  assign _T_197 = _T_195[1]; // @[LZD.scala 39:21]
  assign _T_198 = _T_195[0]; // @[LZD.scala 39:30]
  assign _T_199 = ~ _T_198; // @[LZD.scala 39:27]
  assign _T_200 = _T_197 | _T_199; // @[LZD.scala 39:25]
  assign _T_201 = {_T_196,_T_200}; // @[Cat.scala 29:58]
  assign _T_202 = _T_194[1:0]; // @[LZD.scala 44:32]
  assign _T_203 = _T_202 != 2'h0; // @[LZD.scala 39:14]
  assign _T_204 = _T_202[1]; // @[LZD.scala 39:21]
  assign _T_205 = _T_202[0]; // @[LZD.scala 39:30]
  assign _T_206 = ~ _T_205; // @[LZD.scala 39:27]
  assign _T_207 = _T_204 | _T_206; // @[LZD.scala 39:25]
  assign _T_208 = {_T_203,_T_207}; // @[Cat.scala 29:58]
  assign _T_209 = _T_201[1]; // @[Shift.scala 12:21]
  assign _T_210 = _T_208[1]; // @[Shift.scala 12:21]
  assign _T_211 = _T_209 | _T_210; // @[LZD.scala 49:16]
  assign _T_212 = ~ _T_210; // @[LZD.scala 49:27]
  assign _T_213 = _T_209 | _T_212; // @[LZD.scala 49:25]
  assign _T_214 = _T_201[0:0]; // @[LZD.scala 49:47]
  assign _T_215 = _T_208[0:0]; // @[LZD.scala 49:59]
  assign _T_216 = _T_209 ? _T_214 : _T_215; // @[LZD.scala 49:35]
  assign _T_218 = {_T_211,_T_213,_T_216}; // @[Cat.scala 29:58]
  assign _T_219 = _T_193[2]; // @[Shift.scala 12:21]
  assign _T_220 = _T_218[2]; // @[Shift.scala 12:21]
  assign _T_221 = _T_219 | _T_220; // @[LZD.scala 49:16]
  assign _T_222 = ~ _T_220; // @[LZD.scala 49:27]
  assign _T_223 = _T_219 | _T_222; // @[LZD.scala 49:25]
  assign _T_224 = _T_193[1:0]; // @[LZD.scala 49:47]
  assign _T_225 = _T_218[1:0]; // @[LZD.scala 49:59]
  assign _T_226 = _T_219 ? _T_224 : _T_225; // @[LZD.scala 49:35]
  assign _T_228 = {_T_221,_T_223,_T_226}; // @[Cat.scala 29:58]
  assign _T_229 = _T_167[3:0]; // @[LZD.scala 44:32]
  assign _T_230 = _T_229[3:2]; // @[LZD.scala 43:32]
  assign _T_231 = _T_230 != 2'h0; // @[LZD.scala 39:14]
  assign _T_232 = _T_230[1]; // @[LZD.scala 39:21]
  assign _T_233 = _T_230[0]; // @[LZD.scala 39:30]
  assign _T_234 = ~ _T_233; // @[LZD.scala 39:27]
  assign _T_235 = _T_232 | _T_234; // @[LZD.scala 39:25]
  assign _T_236 = {_T_231,_T_235}; // @[Cat.scala 29:58]
  assign _T_237 = _T_229[1:0]; // @[LZD.scala 44:32]
  assign _T_238 = _T_237 != 2'h0; // @[LZD.scala 39:14]
  assign _T_239 = _T_237[1]; // @[LZD.scala 39:21]
  assign _T_240 = _T_237[0]; // @[LZD.scala 39:30]
  assign _T_241 = ~ _T_240; // @[LZD.scala 39:27]
  assign _T_242 = _T_239 | _T_241; // @[LZD.scala 39:25]
  assign _T_243 = {_T_238,_T_242}; // @[Cat.scala 29:58]
  assign _T_244 = _T_236[1]; // @[Shift.scala 12:21]
  assign _T_245 = _T_243[1]; // @[Shift.scala 12:21]
  assign _T_246 = _T_244 | _T_245; // @[LZD.scala 49:16]
  assign _T_247 = ~ _T_245; // @[LZD.scala 49:27]
  assign _T_248 = _T_244 | _T_247; // @[LZD.scala 49:25]
  assign _T_249 = _T_236[0:0]; // @[LZD.scala 49:47]
  assign _T_250 = _T_243[0:0]; // @[LZD.scala 49:59]
  assign _T_251 = _T_244 ? _T_249 : _T_250; // @[LZD.scala 49:35]
  assign _T_253 = {_T_246,_T_248,_T_251}; // @[Cat.scala 29:58]
  assign _T_254 = _T_228[3]; // @[Shift.scala 12:21]
  assign _T_256 = _T_228[2:0]; // @[LZD.scala 55:32]
  assign _T_257 = _T_254 ? _T_256 : _T_253; // @[LZD.scala 55:20]
  assign _T_258 = {_T_254,_T_257}; // @[Cat.scala 29:58]
  assign _T_259 = ~ _T_258; // @[convert.scala 21:22]
  assign _T_260 = io_B[10:0]; // @[convert.scala 22:36]
  assign _T_261 = _T_259 < 4'hb; // @[Shift.scala 16:24]
  assign _T_263 = _T_259[3]; // @[Shift.scala 12:21]
  assign _T_264 = _T_260[2:0]; // @[Shift.scala 64:52]
  assign _T_266 = {_T_264,8'h0}; // @[Cat.scala 29:58]
  assign _T_267 = _T_263 ? _T_266 : _T_260; // @[Shift.scala 64:27]
  assign _T_268 = _T_259[2:0]; // @[Shift.scala 66:70]
  assign _T_269 = _T_268[2]; // @[Shift.scala 12:21]
  assign _T_270 = _T_267[6:0]; // @[Shift.scala 64:52]
  assign _T_272 = {_T_270,4'h0}; // @[Cat.scala 29:58]
  assign _T_273 = _T_269 ? _T_272 : _T_267; // @[Shift.scala 64:27]
  assign _T_274 = _T_268[1:0]; // @[Shift.scala 66:70]
  assign _T_275 = _T_274[1]; // @[Shift.scala 12:21]
  assign _T_276 = _T_273[8:0]; // @[Shift.scala 64:52]
  assign _T_278 = {_T_276,2'h0}; // @[Cat.scala 29:58]
  assign _T_279 = _T_275 ? _T_278 : _T_273; // @[Shift.scala 64:27]
  assign _T_280 = _T_274[0:0]; // @[Shift.scala 66:70]
  assign _T_282 = _T_279[9:0]; // @[Shift.scala 64:52]
  assign _T_283 = {_T_282,1'h0}; // @[Cat.scala 29:58]
  assign _T_284 = _T_280 ? _T_283 : _T_279; // @[Shift.scala 64:27]
  assign _T_285 = _T_261 ? _T_284 : 11'h0; // @[Shift.scala 16:10]
  assign _T_286 = _T_285[10:10]; // @[convert.scala 23:34]
  assign decB_fraction = _T_285[9:0]; // @[convert.scala 24:34]
  assign _T_288 = _T_164 == 1'h0; // @[convert.scala 25:26]
  assign _T_290 = _T_164 ? _T_259 : _T_258; // @[convert.scala 25:42]
  assign _T_293 = ~ _T_286; // @[convert.scala 26:67]
  assign _T_294 = _T_162 ? _T_293 : _T_286; // @[convert.scala 26:51]
  assign _T_295 = {_T_288,_T_290,_T_294}; // @[Cat.scala 29:58]
  assign _T_297 = io_B[12:0]; // @[convert.scala 29:56]
  assign _T_298 = _T_297 != 13'h0; // @[convert.scala 29:60]
  assign _T_299 = ~ _T_298; // @[convert.scala 29:41]
  assign decB_isNaR = _T_162 & _T_299; // @[convert.scala 29:39]
  assign _T_302 = _T_162 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_302 & _T_299; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_295); // @[convert.scala 32:24]
  assign _T_311 = realC[13]; // @[convert.scala 18:24]
  assign _T_312 = realC[12]; // @[convert.scala 18:40]
  assign _T_313 = _T_311 ^ _T_312; // @[convert.scala 18:36]
  assign _T_314 = realC[12:1]; // @[convert.scala 19:24]
  assign _T_315 = realC[11:0]; // @[convert.scala 19:43]
  assign _T_316 = _T_314 ^ _T_315; // @[convert.scala 19:39]
  assign _T_317 = _T_316[11:4]; // @[LZD.scala 43:32]
  assign _T_318 = _T_317[7:4]; // @[LZD.scala 43:32]
  assign _T_319 = _T_318[3:2]; // @[LZD.scala 43:32]
  assign _T_320 = _T_319 != 2'h0; // @[LZD.scala 39:14]
  assign _T_321 = _T_319[1]; // @[LZD.scala 39:21]
  assign _T_322 = _T_319[0]; // @[LZD.scala 39:30]
  assign _T_323 = ~ _T_322; // @[LZD.scala 39:27]
  assign _T_324 = _T_321 | _T_323; // @[LZD.scala 39:25]
  assign _T_325 = {_T_320,_T_324}; // @[Cat.scala 29:58]
  assign _T_326 = _T_318[1:0]; // @[LZD.scala 44:32]
  assign _T_327 = _T_326 != 2'h0; // @[LZD.scala 39:14]
  assign _T_328 = _T_326[1]; // @[LZD.scala 39:21]
  assign _T_329 = _T_326[0]; // @[LZD.scala 39:30]
  assign _T_330 = ~ _T_329; // @[LZD.scala 39:27]
  assign _T_331 = _T_328 | _T_330; // @[LZD.scala 39:25]
  assign _T_332 = {_T_327,_T_331}; // @[Cat.scala 29:58]
  assign _T_333 = _T_325[1]; // @[Shift.scala 12:21]
  assign _T_334 = _T_332[1]; // @[Shift.scala 12:21]
  assign _T_335 = _T_333 | _T_334; // @[LZD.scala 49:16]
  assign _T_336 = ~ _T_334; // @[LZD.scala 49:27]
  assign _T_337 = _T_333 | _T_336; // @[LZD.scala 49:25]
  assign _T_338 = _T_325[0:0]; // @[LZD.scala 49:47]
  assign _T_339 = _T_332[0:0]; // @[LZD.scala 49:59]
  assign _T_340 = _T_333 ? _T_338 : _T_339; // @[LZD.scala 49:35]
  assign _T_342 = {_T_335,_T_337,_T_340}; // @[Cat.scala 29:58]
  assign _T_343 = _T_317[3:0]; // @[LZD.scala 44:32]
  assign _T_344 = _T_343[3:2]; // @[LZD.scala 43:32]
  assign _T_345 = _T_344 != 2'h0; // @[LZD.scala 39:14]
  assign _T_346 = _T_344[1]; // @[LZD.scala 39:21]
  assign _T_347 = _T_344[0]; // @[LZD.scala 39:30]
  assign _T_348 = ~ _T_347; // @[LZD.scala 39:27]
  assign _T_349 = _T_346 | _T_348; // @[LZD.scala 39:25]
  assign _T_350 = {_T_345,_T_349}; // @[Cat.scala 29:58]
  assign _T_351 = _T_343[1:0]; // @[LZD.scala 44:32]
  assign _T_352 = _T_351 != 2'h0; // @[LZD.scala 39:14]
  assign _T_353 = _T_351[1]; // @[LZD.scala 39:21]
  assign _T_354 = _T_351[0]; // @[LZD.scala 39:30]
  assign _T_355 = ~ _T_354; // @[LZD.scala 39:27]
  assign _T_356 = _T_353 | _T_355; // @[LZD.scala 39:25]
  assign _T_357 = {_T_352,_T_356}; // @[Cat.scala 29:58]
  assign _T_358 = _T_350[1]; // @[Shift.scala 12:21]
  assign _T_359 = _T_357[1]; // @[Shift.scala 12:21]
  assign _T_360 = _T_358 | _T_359; // @[LZD.scala 49:16]
  assign _T_361 = ~ _T_359; // @[LZD.scala 49:27]
  assign _T_362 = _T_358 | _T_361; // @[LZD.scala 49:25]
  assign _T_363 = _T_350[0:0]; // @[LZD.scala 49:47]
  assign _T_364 = _T_357[0:0]; // @[LZD.scala 49:59]
  assign _T_365 = _T_358 ? _T_363 : _T_364; // @[LZD.scala 49:35]
  assign _T_367 = {_T_360,_T_362,_T_365}; // @[Cat.scala 29:58]
  assign _T_368 = _T_342[2]; // @[Shift.scala 12:21]
  assign _T_369 = _T_367[2]; // @[Shift.scala 12:21]
  assign _T_370 = _T_368 | _T_369; // @[LZD.scala 49:16]
  assign _T_371 = ~ _T_369; // @[LZD.scala 49:27]
  assign _T_372 = _T_368 | _T_371; // @[LZD.scala 49:25]
  assign _T_373 = _T_342[1:0]; // @[LZD.scala 49:47]
  assign _T_374 = _T_367[1:0]; // @[LZD.scala 49:59]
  assign _T_375 = _T_368 ? _T_373 : _T_374; // @[LZD.scala 49:35]
  assign _T_377 = {_T_370,_T_372,_T_375}; // @[Cat.scala 29:58]
  assign _T_378 = _T_316[3:0]; // @[LZD.scala 44:32]
  assign _T_379 = _T_378[3:2]; // @[LZD.scala 43:32]
  assign _T_380 = _T_379 != 2'h0; // @[LZD.scala 39:14]
  assign _T_381 = _T_379[1]; // @[LZD.scala 39:21]
  assign _T_382 = _T_379[0]; // @[LZD.scala 39:30]
  assign _T_383 = ~ _T_382; // @[LZD.scala 39:27]
  assign _T_384 = _T_381 | _T_383; // @[LZD.scala 39:25]
  assign _T_385 = {_T_380,_T_384}; // @[Cat.scala 29:58]
  assign _T_386 = _T_378[1:0]; // @[LZD.scala 44:32]
  assign _T_387 = _T_386 != 2'h0; // @[LZD.scala 39:14]
  assign _T_388 = _T_386[1]; // @[LZD.scala 39:21]
  assign _T_389 = _T_386[0]; // @[LZD.scala 39:30]
  assign _T_390 = ~ _T_389; // @[LZD.scala 39:27]
  assign _T_391 = _T_388 | _T_390; // @[LZD.scala 39:25]
  assign _T_392 = {_T_387,_T_391}; // @[Cat.scala 29:58]
  assign _T_393 = _T_385[1]; // @[Shift.scala 12:21]
  assign _T_394 = _T_392[1]; // @[Shift.scala 12:21]
  assign _T_395 = _T_393 | _T_394; // @[LZD.scala 49:16]
  assign _T_396 = ~ _T_394; // @[LZD.scala 49:27]
  assign _T_397 = _T_393 | _T_396; // @[LZD.scala 49:25]
  assign _T_398 = _T_385[0:0]; // @[LZD.scala 49:47]
  assign _T_399 = _T_392[0:0]; // @[LZD.scala 49:59]
  assign _T_400 = _T_393 ? _T_398 : _T_399; // @[LZD.scala 49:35]
  assign _T_402 = {_T_395,_T_397,_T_400}; // @[Cat.scala 29:58]
  assign _T_403 = _T_377[3]; // @[Shift.scala 12:21]
  assign _T_405 = _T_377[2:0]; // @[LZD.scala 55:32]
  assign _T_406 = _T_403 ? _T_405 : _T_402; // @[LZD.scala 55:20]
  assign _T_407 = {_T_403,_T_406}; // @[Cat.scala 29:58]
  assign _T_408 = ~ _T_407; // @[convert.scala 21:22]
  assign _T_409 = realC[10:0]; // @[convert.scala 22:36]
  assign _T_410 = _T_408 < 4'hb; // @[Shift.scala 16:24]
  assign _T_412 = _T_408[3]; // @[Shift.scala 12:21]
  assign _T_413 = _T_409[2:0]; // @[Shift.scala 64:52]
  assign _T_415 = {_T_413,8'h0}; // @[Cat.scala 29:58]
  assign _T_416 = _T_412 ? _T_415 : _T_409; // @[Shift.scala 64:27]
  assign _T_417 = _T_408[2:0]; // @[Shift.scala 66:70]
  assign _T_418 = _T_417[2]; // @[Shift.scala 12:21]
  assign _T_419 = _T_416[6:0]; // @[Shift.scala 64:52]
  assign _T_421 = {_T_419,4'h0}; // @[Cat.scala 29:58]
  assign _T_422 = _T_418 ? _T_421 : _T_416; // @[Shift.scala 64:27]
  assign _T_423 = _T_417[1:0]; // @[Shift.scala 66:70]
  assign _T_424 = _T_423[1]; // @[Shift.scala 12:21]
  assign _T_425 = _T_422[8:0]; // @[Shift.scala 64:52]
  assign _T_427 = {_T_425,2'h0}; // @[Cat.scala 29:58]
  assign _T_428 = _T_424 ? _T_427 : _T_422; // @[Shift.scala 64:27]
  assign _T_429 = _T_423[0:0]; // @[Shift.scala 66:70]
  assign _T_431 = _T_428[9:0]; // @[Shift.scala 64:52]
  assign _T_432 = {_T_431,1'h0}; // @[Cat.scala 29:58]
  assign _T_433 = _T_429 ? _T_432 : _T_428; // @[Shift.scala 64:27]
  assign _T_434 = _T_410 ? _T_433 : 11'h0; // @[Shift.scala 16:10]
  assign _T_435 = _T_434[10:10]; // @[convert.scala 23:34]
  assign decC_fraction = _T_434[9:0]; // @[convert.scala 24:34]
  assign _T_437 = _T_313 == 1'h0; // @[convert.scala 25:26]
  assign _T_439 = _T_313 ? _T_408 : _T_407; // @[convert.scala 25:42]
  assign _T_442 = ~ _T_435; // @[convert.scala 26:67]
  assign _T_443 = _T_311 ? _T_442 : _T_435; // @[convert.scala 26:51]
  assign _T_444 = {_T_437,_T_439,_T_443}; // @[Cat.scala 29:58]
  assign _T_446 = realC[12:0]; // @[convert.scala 29:56]
  assign _T_447 = _T_446 != 13'h0; // @[convert.scala 29:60]
  assign _T_448 = ~ _T_447; // @[convert.scala 29:41]
  assign decC_isNaR = _T_311 & _T_448; // @[convert.scala 29:39]
  assign _T_451 = _T_311 == 1'h0; // @[convert.scala 30:19]
  assign decC_isZero = _T_451 & _T_448; // @[convert.scala 30:41]
  assign decC_scale = $signed(_T_444); // @[convert.scala 32:24]
  assign _T_459 = decA_isNaR | decB_isNaR; // @[PositFMA.scala 58:30]
  assign outIsNaR = _T_459 | decC_isNaR; // @[PositFMA.scala 58:44]
  assign _T_460 = ~ _T_13; // @[PositFMA.scala 59:34]
  assign _T_461 = ~ decA_isZero; // @[PositFMA.scala 59:47]
  assign _T_462 = _T_460 & _T_461; // @[PositFMA.scala 59:45]
  assign _T_464 = {_T_13,_T_462,decA_fraction}; // @[Cat.scala 29:58]
  assign sigA = $signed(_T_464); // @[PositFMA.scala 59:76]
  assign _T_465 = ~ _T_162; // @[PositFMA.scala 60:34]
  assign _T_466 = ~ decB_isZero; // @[PositFMA.scala 60:47]
  assign _T_467 = _T_465 & _T_466; // @[PositFMA.scala 60:45]
  assign _T_469 = {_T_162,_T_467,decB_fraction}; // @[Cat.scala 29:58]
  assign sigB = $signed(_T_469); // @[PositFMA.scala 60:76]
  assign _T_470 = $signed(sigA) * $signed(sigB); // @[PositFMA.scala 61:25]
  assign sigP = $unsigned(_T_470); // @[PositFMA.scala 61:33]
  assign head2 = sigP[23:22]; // @[PositFMA.scala 62:28]
  assign _T_471 = head2[1]; // @[PositFMA.scala 63:31]
  assign _T_472 = ~ _T_471; // @[PositFMA.scala 63:25]
  assign _T_473 = head2[0]; // @[PositFMA.scala 63:42]
  assign addTwo = _T_472 & _T_473; // @[PositFMA.scala 63:35]
  assign _T_474 = sigP[23]; // @[PositFMA.scala 65:23]
  assign _T_475 = sigP[21]; // @[PositFMA.scala 65:49]
  assign addOne = _T_474 ^ _T_475; // @[PositFMA.scala 65:43]
  assign _T_476 = {addTwo,addOne}; // @[Cat.scala 29:58]
  assign expBias = {1'b0,$signed(_T_476)}; // @[PositFMA.scala 66:39]
  assign mulSign = sigP[23:23]; // @[PositFMA.scala 67:28]
  assign _T_477 = $signed(decA_scale) + $signed(decB_scale); // @[PositFMA.scala 69:30]
  assign _GEN_12 = {{4{expBias[2]}},expBias}; // @[PositFMA.scala 69:44]
  assign _T_479 = $signed(_T_477) + $signed(_GEN_12); // @[PositFMA.scala 69:44]
  assign mulScale = $signed(_T_479); // @[PositFMA.scala 69:44]
  assign _T_480 = sigP[21:0]; // @[PositFMA.scala 72:29]
  assign _T_481 = sigP[20:0]; // @[PositFMA.scala 73:29]
  assign _T_482 = {_T_481, 1'h0}; // @[PositFMA.scala 73:48]
  assign mulSigTmp = addOne ? _T_480 : _T_482; // @[PositFMA.scala 70:22]
  assign _T_484 = mulSigTmp[21:21]; // @[PositFMA.scala 77:39]
  assign _T_485 = _T_484 | addTwo; // @[PositFMA.scala 77:43]
  assign _T_486 = mulSigTmp[20:0]; // @[PositFMA.scala 78:39]
  assign mulSig = {mulSign,_T_485,_T_486}; // @[Cat.scala 29:58]
  assign _T_512 = ~ addSign_phase2; // @[PositFMA.scala 107:29]
  assign _T_513 = ~ addZero_phase2; // @[PositFMA.scala 107:47]
  assign _T_514 = _T_512 & _T_513; // @[PositFMA.scala 107:45]
  assign extAddSig = {addSign_phase2,_T_514,addFrac_phase2,11'h0}; // @[Cat.scala 29:58]
  assign _GEN_13 = {{1{addScale_phase2[5]}},addScale_phase2}; // @[PositFMA.scala 111:39]
  assign mulGreater = $signed(mulScale_phase2) > $signed(_GEN_13); // @[PositFMA.scala 111:39]
  assign greaterScale = mulGreater ? $signed(mulScale_phase2) : $signed({{1{addScale_phase2[5]}},addScale_phase2}); // @[PositFMA.scala 112:26]
  assign smallerScale = mulGreater ? $signed({{1{addScale_phase2[5]}},addScale_phase2}) : $signed(mulScale_phase2); // @[PositFMA.scala 113:26]
  assign _T_518 = $signed(greaterScale) - $signed(smallerScale); // @[PositFMA.scala 114:36]
  assign scaleDiff = $signed(_T_518); // @[PositFMA.scala 114:36]
  assign greaterSig = mulGreater ? mulSig_phase2 : extAddSig; // @[PositFMA.scala 115:26]
  assign smallerSigTmp = mulGreater ? extAddSig : mulSig_phase2; // @[PositFMA.scala 116:26]
  assign _T_519 = $unsigned(scaleDiff); // @[PositFMA.scala 117:69]
  assign _T_520 = _T_519 < 7'h17; // @[Shift.scala 39:24]
  assign _T_521 = _T_519[4:0]; // @[Shift.scala 40:44]
  assign _T_522 = smallerSigTmp[22:16]; // @[Shift.scala 90:30]
  assign _T_523 = smallerSigTmp[15:0]; // @[Shift.scala 90:48]
  assign _T_524 = _T_523 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_14 = {{6'd0}, _T_524}; // @[Shift.scala 90:39]
  assign _T_525 = _T_522 | _GEN_14; // @[Shift.scala 90:39]
  assign _T_526 = _T_521[4]; // @[Shift.scala 12:21]
  assign _T_527 = smallerSigTmp[22]; // @[Shift.scala 12:21]
  assign _T_529 = _T_527 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_530 = {_T_529,_T_525}; // @[Cat.scala 29:58]
  assign _T_531 = _T_526 ? _T_530 : smallerSigTmp; // @[Shift.scala 91:22]
  assign _T_532 = _T_521[3:0]; // @[Shift.scala 92:77]
  assign _T_533 = _T_531[22:8]; // @[Shift.scala 90:30]
  assign _T_534 = _T_531[7:0]; // @[Shift.scala 90:48]
  assign _T_535 = _T_534 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_15 = {{14'd0}, _T_535}; // @[Shift.scala 90:39]
  assign _T_536 = _T_533 | _GEN_15; // @[Shift.scala 90:39]
  assign _T_537 = _T_532[3]; // @[Shift.scala 12:21]
  assign _T_538 = _T_531[22]; // @[Shift.scala 12:21]
  assign _T_540 = _T_538 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_541 = {_T_540,_T_536}; // @[Cat.scala 29:58]
  assign _T_542 = _T_537 ? _T_541 : _T_531; // @[Shift.scala 91:22]
  assign _T_543 = _T_532[2:0]; // @[Shift.scala 92:77]
  assign _T_544 = _T_542[22:4]; // @[Shift.scala 90:30]
  assign _T_545 = _T_542[3:0]; // @[Shift.scala 90:48]
  assign _T_546 = _T_545 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_16 = {{18'd0}, _T_546}; // @[Shift.scala 90:39]
  assign _T_547 = _T_544 | _GEN_16; // @[Shift.scala 90:39]
  assign _T_548 = _T_543[2]; // @[Shift.scala 12:21]
  assign _T_549 = _T_542[22]; // @[Shift.scala 12:21]
  assign _T_551 = _T_549 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_552 = {_T_551,_T_547}; // @[Cat.scala 29:58]
  assign _T_553 = _T_548 ? _T_552 : _T_542; // @[Shift.scala 91:22]
  assign _T_554 = _T_543[1:0]; // @[Shift.scala 92:77]
  assign _T_555 = _T_553[22:2]; // @[Shift.scala 90:30]
  assign _T_556 = _T_553[1:0]; // @[Shift.scala 90:48]
  assign _T_557 = _T_556 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_17 = {{20'd0}, _T_557}; // @[Shift.scala 90:39]
  assign _T_558 = _T_555 | _GEN_17; // @[Shift.scala 90:39]
  assign _T_559 = _T_554[1]; // @[Shift.scala 12:21]
  assign _T_560 = _T_553[22]; // @[Shift.scala 12:21]
  assign _T_562 = _T_560 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_563 = {_T_562,_T_558}; // @[Cat.scala 29:58]
  assign _T_564 = _T_559 ? _T_563 : _T_553; // @[Shift.scala 91:22]
  assign _T_565 = _T_554[0:0]; // @[Shift.scala 92:77]
  assign _T_566 = _T_564[22:1]; // @[Shift.scala 90:30]
  assign _T_567 = _T_564[0:0]; // @[Shift.scala 90:48]
  assign _GEN_18 = {{21'd0}, _T_567}; // @[Shift.scala 90:39]
  assign _T_569 = _T_566 | _GEN_18; // @[Shift.scala 90:39]
  assign _T_571 = _T_564[22]; // @[Shift.scala 12:21]
  assign _T_572 = {_T_571,_T_569}; // @[Cat.scala 29:58]
  assign _T_573 = _T_565 ? _T_572 : _T_564; // @[Shift.scala 91:22]
  assign _T_576 = _T_527 ? 23'h7fffff : 23'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_520 ? _T_573 : _T_576; // @[Shift.scala 39:10]
  assign rawSumSig = greaterSig + smallerSig; // @[PositFMA.scala 118:34]
  assign _T_577 = mulSig_phase2[22:22]; // @[PositFMA.scala 119:42]
  assign _T_578 = _T_577 ^ addSign_phase2; // @[PositFMA.scala 119:46]
  assign _T_579 = rawSumSig[23:23]; // @[PositFMA.scala 119:79]
  assign sumSign = _T_578 ^ _T_579; // @[PositFMA.scala 119:63]
  assign _T_581 = greaterSig + smallerSig; // @[PositFMA.scala 120:50]
  assign signSumSig = {sumSign,_T_581}; // @[Cat.scala 29:58]
  assign _T_582 = signSumSig[23:1]; // @[PositFMA.scala 124:33]
  assign _T_583 = signSumSig[22:0]; // @[PositFMA.scala 124:68]
  assign sumXor = _T_582 ^ _T_583; // @[PositFMA.scala 124:51]
  assign _T_584 = sumXor[22:7]; // @[LZD.scala 43:32]
  assign _T_585 = _T_584[15:8]; // @[LZD.scala 43:32]
  assign _T_586 = _T_585[7:4]; // @[LZD.scala 43:32]
  assign _T_587 = _T_586[3:2]; // @[LZD.scala 43:32]
  assign _T_588 = _T_587 != 2'h0; // @[LZD.scala 39:14]
  assign _T_589 = _T_587[1]; // @[LZD.scala 39:21]
  assign _T_590 = _T_587[0]; // @[LZD.scala 39:30]
  assign _T_591 = ~ _T_590; // @[LZD.scala 39:27]
  assign _T_592 = _T_589 | _T_591; // @[LZD.scala 39:25]
  assign _T_593 = {_T_588,_T_592}; // @[Cat.scala 29:58]
  assign _T_594 = _T_586[1:0]; // @[LZD.scala 44:32]
  assign _T_595 = _T_594 != 2'h0; // @[LZD.scala 39:14]
  assign _T_596 = _T_594[1]; // @[LZD.scala 39:21]
  assign _T_597 = _T_594[0]; // @[LZD.scala 39:30]
  assign _T_598 = ~ _T_597; // @[LZD.scala 39:27]
  assign _T_599 = _T_596 | _T_598; // @[LZD.scala 39:25]
  assign _T_600 = {_T_595,_T_599}; // @[Cat.scala 29:58]
  assign _T_601 = _T_593[1]; // @[Shift.scala 12:21]
  assign _T_602 = _T_600[1]; // @[Shift.scala 12:21]
  assign _T_603 = _T_601 | _T_602; // @[LZD.scala 49:16]
  assign _T_604 = ~ _T_602; // @[LZD.scala 49:27]
  assign _T_605 = _T_601 | _T_604; // @[LZD.scala 49:25]
  assign _T_606 = _T_593[0:0]; // @[LZD.scala 49:47]
  assign _T_607 = _T_600[0:0]; // @[LZD.scala 49:59]
  assign _T_608 = _T_601 ? _T_606 : _T_607; // @[LZD.scala 49:35]
  assign _T_610 = {_T_603,_T_605,_T_608}; // @[Cat.scala 29:58]
  assign _T_611 = _T_585[3:0]; // @[LZD.scala 44:32]
  assign _T_612 = _T_611[3:2]; // @[LZD.scala 43:32]
  assign _T_613 = _T_612 != 2'h0; // @[LZD.scala 39:14]
  assign _T_614 = _T_612[1]; // @[LZD.scala 39:21]
  assign _T_615 = _T_612[0]; // @[LZD.scala 39:30]
  assign _T_616 = ~ _T_615; // @[LZD.scala 39:27]
  assign _T_617 = _T_614 | _T_616; // @[LZD.scala 39:25]
  assign _T_618 = {_T_613,_T_617}; // @[Cat.scala 29:58]
  assign _T_619 = _T_611[1:0]; // @[LZD.scala 44:32]
  assign _T_620 = _T_619 != 2'h0; // @[LZD.scala 39:14]
  assign _T_621 = _T_619[1]; // @[LZD.scala 39:21]
  assign _T_622 = _T_619[0]; // @[LZD.scala 39:30]
  assign _T_623 = ~ _T_622; // @[LZD.scala 39:27]
  assign _T_624 = _T_621 | _T_623; // @[LZD.scala 39:25]
  assign _T_625 = {_T_620,_T_624}; // @[Cat.scala 29:58]
  assign _T_626 = _T_618[1]; // @[Shift.scala 12:21]
  assign _T_627 = _T_625[1]; // @[Shift.scala 12:21]
  assign _T_628 = _T_626 | _T_627; // @[LZD.scala 49:16]
  assign _T_629 = ~ _T_627; // @[LZD.scala 49:27]
  assign _T_630 = _T_626 | _T_629; // @[LZD.scala 49:25]
  assign _T_631 = _T_618[0:0]; // @[LZD.scala 49:47]
  assign _T_632 = _T_625[0:0]; // @[LZD.scala 49:59]
  assign _T_633 = _T_626 ? _T_631 : _T_632; // @[LZD.scala 49:35]
  assign _T_635 = {_T_628,_T_630,_T_633}; // @[Cat.scala 29:58]
  assign _T_636 = _T_610[2]; // @[Shift.scala 12:21]
  assign _T_637 = _T_635[2]; // @[Shift.scala 12:21]
  assign _T_638 = _T_636 | _T_637; // @[LZD.scala 49:16]
  assign _T_639 = ~ _T_637; // @[LZD.scala 49:27]
  assign _T_640 = _T_636 | _T_639; // @[LZD.scala 49:25]
  assign _T_641 = _T_610[1:0]; // @[LZD.scala 49:47]
  assign _T_642 = _T_635[1:0]; // @[LZD.scala 49:59]
  assign _T_643 = _T_636 ? _T_641 : _T_642; // @[LZD.scala 49:35]
  assign _T_645 = {_T_638,_T_640,_T_643}; // @[Cat.scala 29:58]
  assign _T_646 = _T_584[7:0]; // @[LZD.scala 44:32]
  assign _T_647 = _T_646[7:4]; // @[LZD.scala 43:32]
  assign _T_648 = _T_647[3:2]; // @[LZD.scala 43:32]
  assign _T_649 = _T_648 != 2'h0; // @[LZD.scala 39:14]
  assign _T_650 = _T_648[1]; // @[LZD.scala 39:21]
  assign _T_651 = _T_648[0]; // @[LZD.scala 39:30]
  assign _T_652 = ~ _T_651; // @[LZD.scala 39:27]
  assign _T_653 = _T_650 | _T_652; // @[LZD.scala 39:25]
  assign _T_654 = {_T_649,_T_653}; // @[Cat.scala 29:58]
  assign _T_655 = _T_647[1:0]; // @[LZD.scala 44:32]
  assign _T_656 = _T_655 != 2'h0; // @[LZD.scala 39:14]
  assign _T_657 = _T_655[1]; // @[LZD.scala 39:21]
  assign _T_658 = _T_655[0]; // @[LZD.scala 39:30]
  assign _T_659 = ~ _T_658; // @[LZD.scala 39:27]
  assign _T_660 = _T_657 | _T_659; // @[LZD.scala 39:25]
  assign _T_661 = {_T_656,_T_660}; // @[Cat.scala 29:58]
  assign _T_662 = _T_654[1]; // @[Shift.scala 12:21]
  assign _T_663 = _T_661[1]; // @[Shift.scala 12:21]
  assign _T_664 = _T_662 | _T_663; // @[LZD.scala 49:16]
  assign _T_665 = ~ _T_663; // @[LZD.scala 49:27]
  assign _T_666 = _T_662 | _T_665; // @[LZD.scala 49:25]
  assign _T_667 = _T_654[0:0]; // @[LZD.scala 49:47]
  assign _T_668 = _T_661[0:0]; // @[LZD.scala 49:59]
  assign _T_669 = _T_662 ? _T_667 : _T_668; // @[LZD.scala 49:35]
  assign _T_671 = {_T_664,_T_666,_T_669}; // @[Cat.scala 29:58]
  assign _T_672 = _T_646[3:0]; // @[LZD.scala 44:32]
  assign _T_673 = _T_672[3:2]; // @[LZD.scala 43:32]
  assign _T_674 = _T_673 != 2'h0; // @[LZD.scala 39:14]
  assign _T_675 = _T_673[1]; // @[LZD.scala 39:21]
  assign _T_676 = _T_673[0]; // @[LZD.scala 39:30]
  assign _T_677 = ~ _T_676; // @[LZD.scala 39:27]
  assign _T_678 = _T_675 | _T_677; // @[LZD.scala 39:25]
  assign _T_679 = {_T_674,_T_678}; // @[Cat.scala 29:58]
  assign _T_680 = _T_672[1:0]; // @[LZD.scala 44:32]
  assign _T_681 = _T_680 != 2'h0; // @[LZD.scala 39:14]
  assign _T_682 = _T_680[1]; // @[LZD.scala 39:21]
  assign _T_683 = _T_680[0]; // @[LZD.scala 39:30]
  assign _T_684 = ~ _T_683; // @[LZD.scala 39:27]
  assign _T_685 = _T_682 | _T_684; // @[LZD.scala 39:25]
  assign _T_686 = {_T_681,_T_685}; // @[Cat.scala 29:58]
  assign _T_687 = _T_679[1]; // @[Shift.scala 12:21]
  assign _T_688 = _T_686[1]; // @[Shift.scala 12:21]
  assign _T_689 = _T_687 | _T_688; // @[LZD.scala 49:16]
  assign _T_690 = ~ _T_688; // @[LZD.scala 49:27]
  assign _T_691 = _T_687 | _T_690; // @[LZD.scala 49:25]
  assign _T_692 = _T_679[0:0]; // @[LZD.scala 49:47]
  assign _T_693 = _T_686[0:0]; // @[LZD.scala 49:59]
  assign _T_694 = _T_687 ? _T_692 : _T_693; // @[LZD.scala 49:35]
  assign _T_696 = {_T_689,_T_691,_T_694}; // @[Cat.scala 29:58]
  assign _T_697 = _T_671[2]; // @[Shift.scala 12:21]
  assign _T_698 = _T_696[2]; // @[Shift.scala 12:21]
  assign _T_699 = _T_697 | _T_698; // @[LZD.scala 49:16]
  assign _T_700 = ~ _T_698; // @[LZD.scala 49:27]
  assign _T_701 = _T_697 | _T_700; // @[LZD.scala 49:25]
  assign _T_702 = _T_671[1:0]; // @[LZD.scala 49:47]
  assign _T_703 = _T_696[1:0]; // @[LZD.scala 49:59]
  assign _T_704 = _T_697 ? _T_702 : _T_703; // @[LZD.scala 49:35]
  assign _T_706 = {_T_699,_T_701,_T_704}; // @[Cat.scala 29:58]
  assign _T_707 = _T_645[3]; // @[Shift.scala 12:21]
  assign _T_708 = _T_706[3]; // @[Shift.scala 12:21]
  assign _T_709 = _T_707 | _T_708; // @[LZD.scala 49:16]
  assign _T_710 = ~ _T_708; // @[LZD.scala 49:27]
  assign _T_711 = _T_707 | _T_710; // @[LZD.scala 49:25]
  assign _T_712 = _T_645[2:0]; // @[LZD.scala 49:47]
  assign _T_713 = _T_706[2:0]; // @[LZD.scala 49:59]
  assign _T_714 = _T_707 ? _T_712 : _T_713; // @[LZD.scala 49:35]
  assign _T_716 = {_T_709,_T_711,_T_714}; // @[Cat.scala 29:58]
  assign _T_717 = sumXor[6:0]; // @[LZD.scala 44:32]
  assign _T_718 = _T_717[6:3]; // @[LZD.scala 43:32]
  assign _T_719 = _T_718[3:2]; // @[LZD.scala 43:32]
  assign _T_720 = _T_719 != 2'h0; // @[LZD.scala 39:14]
  assign _T_721 = _T_719[1]; // @[LZD.scala 39:21]
  assign _T_722 = _T_719[0]; // @[LZD.scala 39:30]
  assign _T_723 = ~ _T_722; // @[LZD.scala 39:27]
  assign _T_724 = _T_721 | _T_723; // @[LZD.scala 39:25]
  assign _T_725 = {_T_720,_T_724}; // @[Cat.scala 29:58]
  assign _T_726 = _T_718[1:0]; // @[LZD.scala 44:32]
  assign _T_727 = _T_726 != 2'h0; // @[LZD.scala 39:14]
  assign _T_728 = _T_726[1]; // @[LZD.scala 39:21]
  assign _T_729 = _T_726[0]; // @[LZD.scala 39:30]
  assign _T_730 = ~ _T_729; // @[LZD.scala 39:27]
  assign _T_731 = _T_728 | _T_730; // @[LZD.scala 39:25]
  assign _T_732 = {_T_727,_T_731}; // @[Cat.scala 29:58]
  assign _T_733 = _T_725[1]; // @[Shift.scala 12:21]
  assign _T_734 = _T_732[1]; // @[Shift.scala 12:21]
  assign _T_735 = _T_733 | _T_734; // @[LZD.scala 49:16]
  assign _T_736 = ~ _T_734; // @[LZD.scala 49:27]
  assign _T_737 = _T_733 | _T_736; // @[LZD.scala 49:25]
  assign _T_738 = _T_725[0:0]; // @[LZD.scala 49:47]
  assign _T_739 = _T_732[0:0]; // @[LZD.scala 49:59]
  assign _T_740 = _T_733 ? _T_738 : _T_739; // @[LZD.scala 49:35]
  assign _T_742 = {_T_735,_T_737,_T_740}; // @[Cat.scala 29:58]
  assign _T_743 = _T_717[2:0]; // @[LZD.scala 44:32]
  assign _T_744 = _T_743[2:1]; // @[LZD.scala 43:32]
  assign _T_745 = _T_744 != 2'h0; // @[LZD.scala 39:14]
  assign _T_746 = _T_744[1]; // @[LZD.scala 39:21]
  assign _T_747 = _T_744[0]; // @[LZD.scala 39:30]
  assign _T_748 = ~ _T_747; // @[LZD.scala 39:27]
  assign _T_749 = _T_746 | _T_748; // @[LZD.scala 39:25]
  assign _T_750 = {_T_745,_T_749}; // @[Cat.scala 29:58]
  assign _T_751 = _T_743[0:0]; // @[LZD.scala 44:32]
  assign _T_753 = _T_750[1]; // @[Shift.scala 12:21]
  assign _T_755 = _T_750[0:0]; // @[LZD.scala 55:32]
  assign _T_756 = _T_753 ? _T_755 : _T_751; // @[LZD.scala 55:20]
  assign _T_757 = {_T_753,_T_756}; // @[Cat.scala 29:58]
  assign _T_758 = _T_742[2]; // @[Shift.scala 12:21]
  assign _T_760 = _T_742[1:0]; // @[LZD.scala 55:32]
  assign _T_761 = _T_758 ? _T_760 : _T_757; // @[LZD.scala 55:20]
  assign _T_763 = _T_716[4]; // @[Shift.scala 12:21]
  assign _T_765 = {1'h1,_T_758,_T_761}; // @[Cat.scala 29:58]
  assign _T_766 = _T_716[3:0]; // @[LZD.scala 55:32]
  assign _T_767 = _T_763 ? _T_766 : _T_765; // @[LZD.scala 55:20]
  assign sumLZD = {_T_763,_T_767}; // @[Cat.scala 29:58]
  assign shiftValue = ~ sumLZD; // @[PositFMA.scala 126:24]
  assign _T_768 = signSumSig[21:0]; // @[PositFMA.scala 127:38]
  assign _T_769 = shiftValue < 5'h16; // @[Shift.scala 16:24]
  assign _T_771 = shiftValue[4]; // @[Shift.scala 12:21]
  assign _T_772 = _T_768[5:0]; // @[Shift.scala 64:52]
  assign _T_774 = {_T_772,16'h0}; // @[Cat.scala 29:58]
  assign _T_775 = _T_771 ? _T_774 : _T_768; // @[Shift.scala 64:27]
  assign _T_776 = shiftValue[3:0]; // @[Shift.scala 66:70]
  assign _T_777 = _T_776[3]; // @[Shift.scala 12:21]
  assign _T_778 = _T_775[13:0]; // @[Shift.scala 64:52]
  assign _T_780 = {_T_778,8'h0}; // @[Cat.scala 29:58]
  assign _T_781 = _T_777 ? _T_780 : _T_775; // @[Shift.scala 64:27]
  assign _T_782 = _T_776[2:0]; // @[Shift.scala 66:70]
  assign _T_783 = _T_782[2]; // @[Shift.scala 12:21]
  assign _T_784 = _T_781[17:0]; // @[Shift.scala 64:52]
  assign _T_786 = {_T_784,4'h0}; // @[Cat.scala 29:58]
  assign _T_787 = _T_783 ? _T_786 : _T_781; // @[Shift.scala 64:27]
  assign _T_788 = _T_782[1:0]; // @[Shift.scala 66:70]
  assign _T_789 = _T_788[1]; // @[Shift.scala 12:21]
  assign _T_790 = _T_787[19:0]; // @[Shift.scala 64:52]
  assign _T_792 = {_T_790,2'h0}; // @[Cat.scala 29:58]
  assign _T_793 = _T_789 ? _T_792 : _T_787; // @[Shift.scala 64:27]
  assign _T_794 = _T_788[0:0]; // @[Shift.scala 66:70]
  assign _T_796 = _T_793[20:0]; // @[Shift.scala 64:52]
  assign _T_797 = {_T_796,1'h0}; // @[Cat.scala 29:58]
  assign _T_798 = _T_794 ? _T_797 : _T_793; // @[Shift.scala 64:27]
  assign normalFracTmp = _T_769 ? _T_798 : 22'h0; // @[Shift.scala 16:10]
  assign _T_800 = $signed(greaterScale) + $signed(7'sh2); // @[PositFMA.scala 130:36]
  assign _T_801 = $signed(_T_800); // @[PositFMA.scala 130:36]
  assign _T_802 = {1'h1,_T_763,_T_767}; // @[Cat.scala 29:58]
  assign _T_803 = $signed(_T_802); // @[PositFMA.scala 130:61]
  assign _GEN_19 = {{1{_T_803[5]}},_T_803}; // @[PositFMA.scala 130:42]
  assign _T_805 = $signed(_T_801) + $signed(_GEN_19); // @[PositFMA.scala 130:42]
  assign sumScale = $signed(_T_805); // @[PositFMA.scala 130:42]
  assign sumFrac = normalFracTmp[21:12]; // @[PositFMA.scala 131:41]
  assign grsTmp = normalFracTmp[11:0]; // @[PositFMA.scala 134:41]
  assign _T_806 = grsTmp[11:10]; // @[PositFMA.scala 137:40]
  assign _T_807 = grsTmp[9:0]; // @[PositFMA.scala 137:56]
  assign _T_808 = _T_807 != 10'h0; // @[PositFMA.scala 137:60]
  assign underflow = $signed(sumScale) < $signed(-7'sh19); // @[PositFMA.scala 144:32]
  assign overflow = $signed(sumScale) > $signed(7'sh18); // @[PositFMA.scala 145:32]
  assign _T_809 = signSumSig != 24'h0; // @[PositFMA.scala 154:32]
  assign decF_isZero = ~ _T_809; // @[PositFMA.scala 154:20]
  assign _T_811 = underflow ? $signed(-7'sh19) : $signed(sumScale); // @[Mux.scala 87:16]
  assign _T_812 = overflow ? $signed(7'sh18) : $signed(_T_811); // @[Mux.scala 87:16]
  assign _GEN_20 = _T_812[5:0]; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  assign decF_scale = $signed(_GEN_20); // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  assign _T_813 = decF_scale[0]; // @[convert.scala 46:61]
  assign _T_814 = ~ _T_813; // @[convert.scala 46:52]
  assign _T_816 = sumSign ? _T_814 : _T_813; // @[convert.scala 46:42]
  assign _T_817 = decF_scale[5:1]; // @[convert.scala 48:34]
  assign _T_818 = _T_817[4:4]; // @[convert.scala 49:36]
  assign _T_820 = ~ _T_817; // @[convert.scala 50:36]
  assign _T_821 = $signed(_T_820); // @[convert.scala 50:36]
  assign _T_822 = _T_818 ? $signed(_T_821) : $signed(_T_817); // @[convert.scala 50:28]
  assign _T_823 = _T_818 ^ sumSign; // @[convert.scala 51:31]
  assign _T_824 = ~ _T_823; // @[convert.scala 52:43]
  assign _T_828 = {_T_824,_T_823,_T_816,sumFrac,_T_806,_T_808}; // @[Cat.scala 29:58]
  assign _T_829 = $unsigned(_T_822); // @[Shift.scala 39:17]
  assign _T_830 = _T_829 < 5'h10; // @[Shift.scala 39:24]
  assign _T_831 = _T_822[3:0]; // @[Shift.scala 40:44]
  assign _T_832 = _T_828[15:8]; // @[Shift.scala 90:30]
  assign _T_833 = _T_828[7:0]; // @[Shift.scala 90:48]
  assign _T_834 = _T_833 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_21 = {{7'd0}, _T_834}; // @[Shift.scala 90:39]
  assign _T_835 = _T_832 | _GEN_21; // @[Shift.scala 90:39]
  assign _T_836 = _T_831[3]; // @[Shift.scala 12:21]
  assign _T_837 = _T_828[15]; // @[Shift.scala 12:21]
  assign _T_839 = _T_837 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_840 = {_T_839,_T_835}; // @[Cat.scala 29:58]
  assign _T_841 = _T_836 ? _T_840 : _T_828; // @[Shift.scala 91:22]
  assign _T_842 = _T_831[2:0]; // @[Shift.scala 92:77]
  assign _T_843 = _T_841[15:4]; // @[Shift.scala 90:30]
  assign _T_844 = _T_841[3:0]; // @[Shift.scala 90:48]
  assign _T_845 = _T_844 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_22 = {{11'd0}, _T_845}; // @[Shift.scala 90:39]
  assign _T_846 = _T_843 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_847 = _T_842[2]; // @[Shift.scala 12:21]
  assign _T_848 = _T_841[15]; // @[Shift.scala 12:21]
  assign _T_850 = _T_848 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_851 = {_T_850,_T_846}; // @[Cat.scala 29:58]
  assign _T_852 = _T_847 ? _T_851 : _T_841; // @[Shift.scala 91:22]
  assign _T_853 = _T_842[1:0]; // @[Shift.scala 92:77]
  assign _T_854 = _T_852[15:2]; // @[Shift.scala 90:30]
  assign _T_855 = _T_852[1:0]; // @[Shift.scala 90:48]
  assign _T_856 = _T_855 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_23 = {{13'd0}, _T_856}; // @[Shift.scala 90:39]
  assign _T_857 = _T_854 | _GEN_23; // @[Shift.scala 90:39]
  assign _T_858 = _T_853[1]; // @[Shift.scala 12:21]
  assign _T_859 = _T_852[15]; // @[Shift.scala 12:21]
  assign _T_861 = _T_859 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_862 = {_T_861,_T_857}; // @[Cat.scala 29:58]
  assign _T_863 = _T_858 ? _T_862 : _T_852; // @[Shift.scala 91:22]
  assign _T_864 = _T_853[0:0]; // @[Shift.scala 92:77]
  assign _T_865 = _T_863[15:1]; // @[Shift.scala 90:30]
  assign _T_866 = _T_863[0:0]; // @[Shift.scala 90:48]
  assign _GEN_24 = {{14'd0}, _T_866}; // @[Shift.scala 90:39]
  assign _T_868 = _T_865 | _GEN_24; // @[Shift.scala 90:39]
  assign _T_870 = _T_863[15]; // @[Shift.scala 12:21]
  assign _T_871 = {_T_870,_T_868}; // @[Cat.scala 29:58]
  assign _T_872 = _T_864 ? _T_871 : _T_863; // @[Shift.scala 91:22]
  assign _T_875 = _T_837 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_876 = _T_830 ? _T_872 : _T_875; // @[Shift.scala 39:10]
  assign _T_877 = _T_876[3]; // @[convert.scala 55:31]
  assign _T_878 = _T_876[2]; // @[convert.scala 56:31]
  assign _T_879 = _T_876[1]; // @[convert.scala 57:31]
  assign _T_880 = _T_876[0]; // @[convert.scala 58:31]
  assign _T_881 = _T_876[15:3]; // @[convert.scala 59:69]
  assign _T_882 = _T_881 != 13'h0; // @[convert.scala 59:81]
  assign _T_883 = ~ _T_882; // @[convert.scala 59:50]
  assign _T_885 = _T_881 == 13'h1fff; // @[convert.scala 60:81]
  assign _T_886 = _T_877 | _T_879; // @[convert.scala 61:44]
  assign _T_887 = _T_886 | _T_880; // @[convert.scala 61:52]
  assign _T_888 = _T_878 & _T_887; // @[convert.scala 61:36]
  assign _T_889 = ~ _T_885; // @[convert.scala 62:63]
  assign _T_890 = _T_889 & _T_888; // @[convert.scala 62:103]
  assign _T_891 = _T_883 | _T_890; // @[convert.scala 62:60]
  assign _GEN_25 = {{12'd0}, _T_891}; // @[convert.scala 63:56]
  assign _T_894 = _T_881 + _GEN_25; // @[convert.scala 63:56]
  assign _T_895 = {sumSign,_T_894}; // @[Cat.scala 29:58]
  assign io_F = _T_903; // @[PositFMA.scala 174:15]
  assign io_outValid = _T_899; // @[PositFMA.scala 173:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  outIsNaR_phase2 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mulSig_phase2 = _RAND_1[22:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  addFrac_phase2 = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mulScale_phase2 = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addScale_phase2 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addSign_phase2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addZero_phase2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  inValid_phase2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_899 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_903 = _RAND_9[13:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (io_inValid) begin
      outIsNaR_phase2 <= outIsNaR;
    end
    if (io_inValid) begin
      mulSig_phase2 <= mulSig;
    end
    if (io_inValid) begin
      addFrac_phase2 <= decC_fraction;
    end
    if (io_inValid) begin
      mulScale_phase2 <= mulScale;
    end
    if (io_inValid) begin
      addScale_phase2 <= decC_scale;
    end
    if (io_inValid) begin
      addSign_phase2 <= _T_311;
    end
    if (io_inValid) begin
      addZero_phase2 <= decC_isZero;
    end
    if (reset) begin
      inValid_phase2 <= 1'h0;
    end else begin
      inValid_phase2 <= io_inValid;
    end
    if (reset) begin
      _T_899 <= 1'h0;
    end else begin
      _T_899 <= inValid_phase2;
    end
    if (inValid_phase2) begin
      if (outIsNaR_phase2) begin
        _T_903 <= 14'h2000;
      end else begin
        if (decF_isZero) begin
          _T_903 <= 14'h0;
        end else begin
          _T_903 <= _T_895;
        end
      end
    end
  end
endmodule
