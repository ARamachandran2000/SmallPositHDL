module PositFMA30_3(
  input         clock,
  input         reset,
  input         io_inValid,
  input  [1:0]  io_fmaOp,
  input  [29:0] io_A,
  input  [29:0] io_B,
  input  [29:0] io_C,
  output [29:0] io_F,
  output        io_outValid
);
  wire  _T; // @[PositFMA.scala 47:36]
  wire [29:0] _T_2; // @[Bitwise.scala 71:12]
  wire [29:0] _T_3; // @[PositFMA.scala 47:41]
  wire [29:0] _GEN_10; // @[PositFMA.scala 47:49]
  wire [29:0] realA; // @[PositFMA.scala 47:49]
  wire  _T_6; // @[PositFMA.scala 48:36]
  wire [29:0] _T_8; // @[Bitwise.scala 71:12]
  wire [29:0] _T_9; // @[PositFMA.scala 48:41]
  wire [29:0] _GEN_11; // @[PositFMA.scala 48:49]
  wire [29:0] realC; // @[PositFMA.scala 48:49]
  wire  _T_13; // @[convert.scala 18:24]
  wire  _T_14; // @[convert.scala 18:40]
  wire  _T_15; // @[convert.scala 18:36]
  wire [27:0] _T_16; // @[convert.scala 19:24]
  wire [27:0] _T_17; // @[convert.scala 19:43]
  wire [27:0] _T_18; // @[convert.scala 19:39]
  wire [15:0] _T_19; // @[LZD.scala 43:32]
  wire [7:0] _T_20; // @[LZD.scala 43:32]
  wire [3:0] _T_21; // @[LZD.scala 43:32]
  wire [1:0] _T_22; // @[LZD.scala 43:32]
  wire  _T_23; // @[LZD.scala 39:14]
  wire  _T_24; // @[LZD.scala 39:21]
  wire  _T_25; // @[LZD.scala 39:30]
  wire  _T_26; // @[LZD.scala 39:27]
  wire  _T_27; // @[LZD.scala 39:25]
  wire [1:0] _T_28; // @[Cat.scala 29:58]
  wire [1:0] _T_29; // @[LZD.scala 44:32]
  wire  _T_30; // @[LZD.scala 39:14]
  wire  _T_31; // @[LZD.scala 39:21]
  wire  _T_32; // @[LZD.scala 39:30]
  wire  _T_33; // @[LZD.scala 39:27]
  wire  _T_34; // @[LZD.scala 39:25]
  wire [1:0] _T_35; // @[Cat.scala 29:58]
  wire  _T_36; // @[Shift.scala 12:21]
  wire  _T_37; // @[Shift.scala 12:21]
  wire  _T_38; // @[LZD.scala 49:16]
  wire  _T_39; // @[LZD.scala 49:27]
  wire  _T_40; // @[LZD.scala 49:25]
  wire  _T_41; // @[LZD.scala 49:47]
  wire  _T_42; // @[LZD.scala 49:59]
  wire  _T_43; // @[LZD.scala 49:35]
  wire [2:0] _T_45; // @[Cat.scala 29:58]
  wire [3:0] _T_46; // @[LZD.scala 44:32]
  wire [1:0] _T_47; // @[LZD.scala 43:32]
  wire  _T_48; // @[LZD.scala 39:14]
  wire  _T_49; // @[LZD.scala 39:21]
  wire  _T_50; // @[LZD.scala 39:30]
  wire  _T_51; // @[LZD.scala 39:27]
  wire  _T_52; // @[LZD.scala 39:25]
  wire [1:0] _T_53; // @[Cat.scala 29:58]
  wire [1:0] _T_54; // @[LZD.scala 44:32]
  wire  _T_55; // @[LZD.scala 39:14]
  wire  _T_56; // @[LZD.scala 39:21]
  wire  _T_57; // @[LZD.scala 39:30]
  wire  _T_58; // @[LZD.scala 39:27]
  wire  _T_59; // @[LZD.scala 39:25]
  wire [1:0] _T_60; // @[Cat.scala 29:58]
  wire  _T_61; // @[Shift.scala 12:21]
  wire  _T_62; // @[Shift.scala 12:21]
  wire  _T_63; // @[LZD.scala 49:16]
  wire  _T_64; // @[LZD.scala 49:27]
  wire  _T_65; // @[LZD.scala 49:25]
  wire  _T_66; // @[LZD.scala 49:47]
  wire  _T_67; // @[LZD.scala 49:59]
  wire  _T_68; // @[LZD.scala 49:35]
  wire [2:0] _T_70; // @[Cat.scala 29:58]
  wire  _T_71; // @[Shift.scala 12:21]
  wire  _T_72; // @[Shift.scala 12:21]
  wire  _T_73; // @[LZD.scala 49:16]
  wire  _T_74; // @[LZD.scala 49:27]
  wire  _T_75; // @[LZD.scala 49:25]
  wire [1:0] _T_76; // @[LZD.scala 49:47]
  wire [1:0] _T_77; // @[LZD.scala 49:59]
  wire [1:0] _T_78; // @[LZD.scala 49:35]
  wire [3:0] _T_80; // @[Cat.scala 29:58]
  wire [7:0] _T_81; // @[LZD.scala 44:32]
  wire [3:0] _T_82; // @[LZD.scala 43:32]
  wire [1:0] _T_83; // @[LZD.scala 43:32]
  wire  _T_84; // @[LZD.scala 39:14]
  wire  _T_85; // @[LZD.scala 39:21]
  wire  _T_86; // @[LZD.scala 39:30]
  wire  _T_87; // @[LZD.scala 39:27]
  wire  _T_88; // @[LZD.scala 39:25]
  wire [1:0] _T_89; // @[Cat.scala 29:58]
  wire [1:0] _T_90; // @[LZD.scala 44:32]
  wire  _T_91; // @[LZD.scala 39:14]
  wire  _T_92; // @[LZD.scala 39:21]
  wire  _T_93; // @[LZD.scala 39:30]
  wire  _T_94; // @[LZD.scala 39:27]
  wire  _T_95; // @[LZD.scala 39:25]
  wire [1:0] _T_96; // @[Cat.scala 29:58]
  wire  _T_97; // @[Shift.scala 12:21]
  wire  _T_98; // @[Shift.scala 12:21]
  wire  _T_99; // @[LZD.scala 49:16]
  wire  _T_100; // @[LZD.scala 49:27]
  wire  _T_101; // @[LZD.scala 49:25]
  wire  _T_102; // @[LZD.scala 49:47]
  wire  _T_103; // @[LZD.scala 49:59]
  wire  _T_104; // @[LZD.scala 49:35]
  wire [2:0] _T_106; // @[Cat.scala 29:58]
  wire [3:0] _T_107; // @[LZD.scala 44:32]
  wire [1:0] _T_108; // @[LZD.scala 43:32]
  wire  _T_109; // @[LZD.scala 39:14]
  wire  _T_110; // @[LZD.scala 39:21]
  wire  _T_111; // @[LZD.scala 39:30]
  wire  _T_112; // @[LZD.scala 39:27]
  wire  _T_113; // @[LZD.scala 39:25]
  wire [1:0] _T_114; // @[Cat.scala 29:58]
  wire [1:0] _T_115; // @[LZD.scala 44:32]
  wire  _T_116; // @[LZD.scala 39:14]
  wire  _T_117; // @[LZD.scala 39:21]
  wire  _T_118; // @[LZD.scala 39:30]
  wire  _T_119; // @[LZD.scala 39:27]
  wire  _T_120; // @[LZD.scala 39:25]
  wire [1:0] _T_121; // @[Cat.scala 29:58]
  wire  _T_122; // @[Shift.scala 12:21]
  wire  _T_123; // @[Shift.scala 12:21]
  wire  _T_124; // @[LZD.scala 49:16]
  wire  _T_125; // @[LZD.scala 49:27]
  wire  _T_126; // @[LZD.scala 49:25]
  wire  _T_127; // @[LZD.scala 49:47]
  wire  _T_128; // @[LZD.scala 49:59]
  wire  _T_129; // @[LZD.scala 49:35]
  wire [2:0] _T_131; // @[Cat.scala 29:58]
  wire  _T_132; // @[Shift.scala 12:21]
  wire  _T_133; // @[Shift.scala 12:21]
  wire  _T_134; // @[LZD.scala 49:16]
  wire  _T_135; // @[LZD.scala 49:27]
  wire  _T_136; // @[LZD.scala 49:25]
  wire [1:0] _T_137; // @[LZD.scala 49:47]
  wire [1:0] _T_138; // @[LZD.scala 49:59]
  wire [1:0] _T_139; // @[LZD.scala 49:35]
  wire [3:0] _T_141; // @[Cat.scala 29:58]
  wire  _T_142; // @[Shift.scala 12:21]
  wire  _T_143; // @[Shift.scala 12:21]
  wire  _T_144; // @[LZD.scala 49:16]
  wire  _T_145; // @[LZD.scala 49:27]
  wire  _T_146; // @[LZD.scala 49:25]
  wire [2:0] _T_147; // @[LZD.scala 49:47]
  wire [2:0] _T_148; // @[LZD.scala 49:59]
  wire [2:0] _T_149; // @[LZD.scala 49:35]
  wire [4:0] _T_151; // @[Cat.scala 29:58]
  wire [11:0] _T_152; // @[LZD.scala 44:32]
  wire [7:0] _T_153; // @[LZD.scala 43:32]
  wire [3:0] _T_154; // @[LZD.scala 43:32]
  wire [1:0] _T_155; // @[LZD.scala 43:32]
  wire  _T_156; // @[LZD.scala 39:14]
  wire  _T_157; // @[LZD.scala 39:21]
  wire  _T_158; // @[LZD.scala 39:30]
  wire  _T_159; // @[LZD.scala 39:27]
  wire  _T_160; // @[LZD.scala 39:25]
  wire [1:0] _T_161; // @[Cat.scala 29:58]
  wire [1:0] _T_162; // @[LZD.scala 44:32]
  wire  _T_163; // @[LZD.scala 39:14]
  wire  _T_164; // @[LZD.scala 39:21]
  wire  _T_165; // @[LZD.scala 39:30]
  wire  _T_166; // @[LZD.scala 39:27]
  wire  _T_167; // @[LZD.scala 39:25]
  wire [1:0] _T_168; // @[Cat.scala 29:58]
  wire  _T_169; // @[Shift.scala 12:21]
  wire  _T_170; // @[Shift.scala 12:21]
  wire  _T_171; // @[LZD.scala 49:16]
  wire  _T_172; // @[LZD.scala 49:27]
  wire  _T_173; // @[LZD.scala 49:25]
  wire  _T_174; // @[LZD.scala 49:47]
  wire  _T_175; // @[LZD.scala 49:59]
  wire  _T_176; // @[LZD.scala 49:35]
  wire [2:0] _T_178; // @[Cat.scala 29:58]
  wire [3:0] _T_179; // @[LZD.scala 44:32]
  wire [1:0] _T_180; // @[LZD.scala 43:32]
  wire  _T_181; // @[LZD.scala 39:14]
  wire  _T_182; // @[LZD.scala 39:21]
  wire  _T_183; // @[LZD.scala 39:30]
  wire  _T_184; // @[LZD.scala 39:27]
  wire  _T_185; // @[LZD.scala 39:25]
  wire [1:0] _T_186; // @[Cat.scala 29:58]
  wire [1:0] _T_187; // @[LZD.scala 44:32]
  wire  _T_188; // @[LZD.scala 39:14]
  wire  _T_189; // @[LZD.scala 39:21]
  wire  _T_190; // @[LZD.scala 39:30]
  wire  _T_191; // @[LZD.scala 39:27]
  wire  _T_192; // @[LZD.scala 39:25]
  wire [1:0] _T_193; // @[Cat.scala 29:58]
  wire  _T_194; // @[Shift.scala 12:21]
  wire  _T_195; // @[Shift.scala 12:21]
  wire  _T_196; // @[LZD.scala 49:16]
  wire  _T_197; // @[LZD.scala 49:27]
  wire  _T_198; // @[LZD.scala 49:25]
  wire  _T_199; // @[LZD.scala 49:47]
  wire  _T_200; // @[LZD.scala 49:59]
  wire  _T_201; // @[LZD.scala 49:35]
  wire [2:0] _T_203; // @[Cat.scala 29:58]
  wire  _T_204; // @[Shift.scala 12:21]
  wire  _T_205; // @[Shift.scala 12:21]
  wire  _T_206; // @[LZD.scala 49:16]
  wire  _T_207; // @[LZD.scala 49:27]
  wire  _T_208; // @[LZD.scala 49:25]
  wire [1:0] _T_209; // @[LZD.scala 49:47]
  wire [1:0] _T_210; // @[LZD.scala 49:59]
  wire [1:0] _T_211; // @[LZD.scala 49:35]
  wire [3:0] _T_213; // @[Cat.scala 29:58]
  wire [3:0] _T_214; // @[LZD.scala 44:32]
  wire [1:0] _T_215; // @[LZD.scala 43:32]
  wire  _T_216; // @[LZD.scala 39:14]
  wire  _T_217; // @[LZD.scala 39:21]
  wire  _T_218; // @[LZD.scala 39:30]
  wire  _T_219; // @[LZD.scala 39:27]
  wire  _T_220; // @[LZD.scala 39:25]
  wire [1:0] _T_221; // @[Cat.scala 29:58]
  wire [1:0] _T_222; // @[LZD.scala 44:32]
  wire  _T_223; // @[LZD.scala 39:14]
  wire  _T_224; // @[LZD.scala 39:21]
  wire  _T_225; // @[LZD.scala 39:30]
  wire  _T_226; // @[LZD.scala 39:27]
  wire  _T_227; // @[LZD.scala 39:25]
  wire [1:0] _T_228; // @[Cat.scala 29:58]
  wire  _T_229; // @[Shift.scala 12:21]
  wire  _T_230; // @[Shift.scala 12:21]
  wire  _T_231; // @[LZD.scala 49:16]
  wire  _T_232; // @[LZD.scala 49:27]
  wire  _T_233; // @[LZD.scala 49:25]
  wire  _T_234; // @[LZD.scala 49:47]
  wire  _T_235; // @[LZD.scala 49:59]
  wire  _T_236; // @[LZD.scala 49:35]
  wire [2:0] _T_238; // @[Cat.scala 29:58]
  wire  _T_239; // @[Shift.scala 12:21]
  wire [2:0] _T_241; // @[LZD.scala 55:32]
  wire [2:0] _T_242; // @[LZD.scala 55:20]
  wire [3:0] _T_243; // @[Cat.scala 29:58]
  wire  _T_244; // @[Shift.scala 12:21]
  wire [3:0] _T_246; // @[LZD.scala 55:32]
  wire [3:0] _T_247; // @[LZD.scala 55:20]
  wire [4:0] _T_248; // @[Cat.scala 29:58]
  wire [4:0] _T_249; // @[convert.scala 21:22]
  wire [26:0] _T_250; // @[convert.scala 22:36]
  wire  _T_251; // @[Shift.scala 16:24]
  wire  _T_253; // @[Shift.scala 12:21]
  wire [10:0] _T_254; // @[Shift.scala 64:52]
  wire [26:0] _T_256; // @[Cat.scala 29:58]
  wire [26:0] _T_257; // @[Shift.scala 64:27]
  wire [3:0] _T_258; // @[Shift.scala 66:70]
  wire  _T_259; // @[Shift.scala 12:21]
  wire [18:0] _T_260; // @[Shift.scala 64:52]
  wire [26:0] _T_262; // @[Cat.scala 29:58]
  wire [26:0] _T_263; // @[Shift.scala 64:27]
  wire [2:0] _T_264; // @[Shift.scala 66:70]
  wire  _T_265; // @[Shift.scala 12:21]
  wire [22:0] _T_266; // @[Shift.scala 64:52]
  wire [26:0] _T_268; // @[Cat.scala 29:58]
  wire [26:0] _T_269; // @[Shift.scala 64:27]
  wire [1:0] _T_270; // @[Shift.scala 66:70]
  wire  _T_271; // @[Shift.scala 12:21]
  wire [24:0] _T_272; // @[Shift.scala 64:52]
  wire [26:0] _T_274; // @[Cat.scala 29:58]
  wire [26:0] _T_275; // @[Shift.scala 64:27]
  wire  _T_276; // @[Shift.scala 66:70]
  wire [25:0] _T_278; // @[Shift.scala 64:52]
  wire [26:0] _T_279; // @[Cat.scala 29:58]
  wire [26:0] _T_280; // @[Shift.scala 64:27]
  wire [26:0] _T_281; // @[Shift.scala 16:10]
  wire [2:0] _T_282; // @[convert.scala 23:34]
  wire [23:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_284; // @[convert.scala 25:26]
  wire [4:0] _T_286; // @[convert.scala 25:42]
  wire [2:0] _T_289; // @[convert.scala 26:67]
  wire [2:0] _T_290; // @[convert.scala 26:51]
  wire [8:0] _T_291; // @[Cat.scala 29:58]
  wire [28:0] _T_293; // @[convert.scala 29:56]
  wire  _T_294; // @[convert.scala 29:60]
  wire  _T_295; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_298; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [8:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_307; // @[convert.scala 18:24]
  wire  _T_308; // @[convert.scala 18:40]
  wire  _T_309; // @[convert.scala 18:36]
  wire [27:0] _T_310; // @[convert.scala 19:24]
  wire [27:0] _T_311; // @[convert.scala 19:43]
  wire [27:0] _T_312; // @[convert.scala 19:39]
  wire [15:0] _T_313; // @[LZD.scala 43:32]
  wire [7:0] _T_314; // @[LZD.scala 43:32]
  wire [3:0] _T_315; // @[LZD.scala 43:32]
  wire [1:0] _T_316; // @[LZD.scala 43:32]
  wire  _T_317; // @[LZD.scala 39:14]
  wire  _T_318; // @[LZD.scala 39:21]
  wire  _T_319; // @[LZD.scala 39:30]
  wire  _T_320; // @[LZD.scala 39:27]
  wire  _T_321; // @[LZD.scala 39:25]
  wire [1:0] _T_322; // @[Cat.scala 29:58]
  wire [1:0] _T_323; // @[LZD.scala 44:32]
  wire  _T_324; // @[LZD.scala 39:14]
  wire  _T_325; // @[LZD.scala 39:21]
  wire  _T_326; // @[LZD.scala 39:30]
  wire  _T_327; // @[LZD.scala 39:27]
  wire  _T_328; // @[LZD.scala 39:25]
  wire [1:0] _T_329; // @[Cat.scala 29:58]
  wire  _T_330; // @[Shift.scala 12:21]
  wire  _T_331; // @[Shift.scala 12:21]
  wire  _T_332; // @[LZD.scala 49:16]
  wire  _T_333; // @[LZD.scala 49:27]
  wire  _T_334; // @[LZD.scala 49:25]
  wire  _T_335; // @[LZD.scala 49:47]
  wire  _T_336; // @[LZD.scala 49:59]
  wire  _T_337; // @[LZD.scala 49:35]
  wire [2:0] _T_339; // @[Cat.scala 29:58]
  wire [3:0] _T_340; // @[LZD.scala 44:32]
  wire [1:0] _T_341; // @[LZD.scala 43:32]
  wire  _T_342; // @[LZD.scala 39:14]
  wire  _T_343; // @[LZD.scala 39:21]
  wire  _T_344; // @[LZD.scala 39:30]
  wire  _T_345; // @[LZD.scala 39:27]
  wire  _T_346; // @[LZD.scala 39:25]
  wire [1:0] _T_347; // @[Cat.scala 29:58]
  wire [1:0] _T_348; // @[LZD.scala 44:32]
  wire  _T_349; // @[LZD.scala 39:14]
  wire  _T_350; // @[LZD.scala 39:21]
  wire  _T_351; // @[LZD.scala 39:30]
  wire  _T_352; // @[LZD.scala 39:27]
  wire  _T_353; // @[LZD.scala 39:25]
  wire [1:0] _T_354; // @[Cat.scala 29:58]
  wire  _T_355; // @[Shift.scala 12:21]
  wire  _T_356; // @[Shift.scala 12:21]
  wire  _T_357; // @[LZD.scala 49:16]
  wire  _T_358; // @[LZD.scala 49:27]
  wire  _T_359; // @[LZD.scala 49:25]
  wire  _T_360; // @[LZD.scala 49:47]
  wire  _T_361; // @[LZD.scala 49:59]
  wire  _T_362; // @[LZD.scala 49:35]
  wire [2:0] _T_364; // @[Cat.scala 29:58]
  wire  _T_365; // @[Shift.scala 12:21]
  wire  _T_366; // @[Shift.scala 12:21]
  wire  _T_367; // @[LZD.scala 49:16]
  wire  _T_368; // @[LZD.scala 49:27]
  wire  _T_369; // @[LZD.scala 49:25]
  wire [1:0] _T_370; // @[LZD.scala 49:47]
  wire [1:0] _T_371; // @[LZD.scala 49:59]
  wire [1:0] _T_372; // @[LZD.scala 49:35]
  wire [3:0] _T_374; // @[Cat.scala 29:58]
  wire [7:0] _T_375; // @[LZD.scala 44:32]
  wire [3:0] _T_376; // @[LZD.scala 43:32]
  wire [1:0] _T_377; // @[LZD.scala 43:32]
  wire  _T_378; // @[LZD.scala 39:14]
  wire  _T_379; // @[LZD.scala 39:21]
  wire  _T_380; // @[LZD.scala 39:30]
  wire  _T_381; // @[LZD.scala 39:27]
  wire  _T_382; // @[LZD.scala 39:25]
  wire [1:0] _T_383; // @[Cat.scala 29:58]
  wire [1:0] _T_384; // @[LZD.scala 44:32]
  wire  _T_385; // @[LZD.scala 39:14]
  wire  _T_386; // @[LZD.scala 39:21]
  wire  _T_387; // @[LZD.scala 39:30]
  wire  _T_388; // @[LZD.scala 39:27]
  wire  _T_389; // @[LZD.scala 39:25]
  wire [1:0] _T_390; // @[Cat.scala 29:58]
  wire  _T_391; // @[Shift.scala 12:21]
  wire  _T_392; // @[Shift.scala 12:21]
  wire  _T_393; // @[LZD.scala 49:16]
  wire  _T_394; // @[LZD.scala 49:27]
  wire  _T_395; // @[LZD.scala 49:25]
  wire  _T_396; // @[LZD.scala 49:47]
  wire  _T_397; // @[LZD.scala 49:59]
  wire  _T_398; // @[LZD.scala 49:35]
  wire [2:0] _T_400; // @[Cat.scala 29:58]
  wire [3:0] _T_401; // @[LZD.scala 44:32]
  wire [1:0] _T_402; // @[LZD.scala 43:32]
  wire  _T_403; // @[LZD.scala 39:14]
  wire  _T_404; // @[LZD.scala 39:21]
  wire  _T_405; // @[LZD.scala 39:30]
  wire  _T_406; // @[LZD.scala 39:27]
  wire  _T_407; // @[LZD.scala 39:25]
  wire [1:0] _T_408; // @[Cat.scala 29:58]
  wire [1:0] _T_409; // @[LZD.scala 44:32]
  wire  _T_410; // @[LZD.scala 39:14]
  wire  _T_411; // @[LZD.scala 39:21]
  wire  _T_412; // @[LZD.scala 39:30]
  wire  _T_413; // @[LZD.scala 39:27]
  wire  _T_414; // @[LZD.scala 39:25]
  wire [1:0] _T_415; // @[Cat.scala 29:58]
  wire  _T_416; // @[Shift.scala 12:21]
  wire  _T_417; // @[Shift.scala 12:21]
  wire  _T_418; // @[LZD.scala 49:16]
  wire  _T_419; // @[LZD.scala 49:27]
  wire  _T_420; // @[LZD.scala 49:25]
  wire  _T_421; // @[LZD.scala 49:47]
  wire  _T_422; // @[LZD.scala 49:59]
  wire  _T_423; // @[LZD.scala 49:35]
  wire [2:0] _T_425; // @[Cat.scala 29:58]
  wire  _T_426; // @[Shift.scala 12:21]
  wire  _T_427; // @[Shift.scala 12:21]
  wire  _T_428; // @[LZD.scala 49:16]
  wire  _T_429; // @[LZD.scala 49:27]
  wire  _T_430; // @[LZD.scala 49:25]
  wire [1:0] _T_431; // @[LZD.scala 49:47]
  wire [1:0] _T_432; // @[LZD.scala 49:59]
  wire [1:0] _T_433; // @[LZD.scala 49:35]
  wire [3:0] _T_435; // @[Cat.scala 29:58]
  wire  _T_436; // @[Shift.scala 12:21]
  wire  _T_437; // @[Shift.scala 12:21]
  wire  _T_438; // @[LZD.scala 49:16]
  wire  _T_439; // @[LZD.scala 49:27]
  wire  _T_440; // @[LZD.scala 49:25]
  wire [2:0] _T_441; // @[LZD.scala 49:47]
  wire [2:0] _T_442; // @[LZD.scala 49:59]
  wire [2:0] _T_443; // @[LZD.scala 49:35]
  wire [4:0] _T_445; // @[Cat.scala 29:58]
  wire [11:0] _T_446; // @[LZD.scala 44:32]
  wire [7:0] _T_447; // @[LZD.scala 43:32]
  wire [3:0] _T_448; // @[LZD.scala 43:32]
  wire [1:0] _T_449; // @[LZD.scala 43:32]
  wire  _T_450; // @[LZD.scala 39:14]
  wire  _T_451; // @[LZD.scala 39:21]
  wire  _T_452; // @[LZD.scala 39:30]
  wire  _T_453; // @[LZD.scala 39:27]
  wire  _T_454; // @[LZD.scala 39:25]
  wire [1:0] _T_455; // @[Cat.scala 29:58]
  wire [1:0] _T_456; // @[LZD.scala 44:32]
  wire  _T_457; // @[LZD.scala 39:14]
  wire  _T_458; // @[LZD.scala 39:21]
  wire  _T_459; // @[LZD.scala 39:30]
  wire  _T_460; // @[LZD.scala 39:27]
  wire  _T_461; // @[LZD.scala 39:25]
  wire [1:0] _T_462; // @[Cat.scala 29:58]
  wire  _T_463; // @[Shift.scala 12:21]
  wire  _T_464; // @[Shift.scala 12:21]
  wire  _T_465; // @[LZD.scala 49:16]
  wire  _T_466; // @[LZD.scala 49:27]
  wire  _T_467; // @[LZD.scala 49:25]
  wire  _T_468; // @[LZD.scala 49:47]
  wire  _T_469; // @[LZD.scala 49:59]
  wire  _T_470; // @[LZD.scala 49:35]
  wire [2:0] _T_472; // @[Cat.scala 29:58]
  wire [3:0] _T_473; // @[LZD.scala 44:32]
  wire [1:0] _T_474; // @[LZD.scala 43:32]
  wire  _T_475; // @[LZD.scala 39:14]
  wire  _T_476; // @[LZD.scala 39:21]
  wire  _T_477; // @[LZD.scala 39:30]
  wire  _T_478; // @[LZD.scala 39:27]
  wire  _T_479; // @[LZD.scala 39:25]
  wire [1:0] _T_480; // @[Cat.scala 29:58]
  wire [1:0] _T_481; // @[LZD.scala 44:32]
  wire  _T_482; // @[LZD.scala 39:14]
  wire  _T_483; // @[LZD.scala 39:21]
  wire  _T_484; // @[LZD.scala 39:30]
  wire  _T_485; // @[LZD.scala 39:27]
  wire  _T_486; // @[LZD.scala 39:25]
  wire [1:0] _T_487; // @[Cat.scala 29:58]
  wire  _T_488; // @[Shift.scala 12:21]
  wire  _T_489; // @[Shift.scala 12:21]
  wire  _T_490; // @[LZD.scala 49:16]
  wire  _T_491; // @[LZD.scala 49:27]
  wire  _T_492; // @[LZD.scala 49:25]
  wire  _T_493; // @[LZD.scala 49:47]
  wire  _T_494; // @[LZD.scala 49:59]
  wire  _T_495; // @[LZD.scala 49:35]
  wire [2:0] _T_497; // @[Cat.scala 29:58]
  wire  _T_498; // @[Shift.scala 12:21]
  wire  _T_499; // @[Shift.scala 12:21]
  wire  _T_500; // @[LZD.scala 49:16]
  wire  _T_501; // @[LZD.scala 49:27]
  wire  _T_502; // @[LZD.scala 49:25]
  wire [1:0] _T_503; // @[LZD.scala 49:47]
  wire [1:0] _T_504; // @[LZD.scala 49:59]
  wire [1:0] _T_505; // @[LZD.scala 49:35]
  wire [3:0] _T_507; // @[Cat.scala 29:58]
  wire [3:0] _T_508; // @[LZD.scala 44:32]
  wire [1:0] _T_509; // @[LZD.scala 43:32]
  wire  _T_510; // @[LZD.scala 39:14]
  wire  _T_511; // @[LZD.scala 39:21]
  wire  _T_512; // @[LZD.scala 39:30]
  wire  _T_513; // @[LZD.scala 39:27]
  wire  _T_514; // @[LZD.scala 39:25]
  wire [1:0] _T_515; // @[Cat.scala 29:58]
  wire [1:0] _T_516; // @[LZD.scala 44:32]
  wire  _T_517; // @[LZD.scala 39:14]
  wire  _T_518; // @[LZD.scala 39:21]
  wire  _T_519; // @[LZD.scala 39:30]
  wire  _T_520; // @[LZD.scala 39:27]
  wire  _T_521; // @[LZD.scala 39:25]
  wire [1:0] _T_522; // @[Cat.scala 29:58]
  wire  _T_523; // @[Shift.scala 12:21]
  wire  _T_524; // @[Shift.scala 12:21]
  wire  _T_525; // @[LZD.scala 49:16]
  wire  _T_526; // @[LZD.scala 49:27]
  wire  _T_527; // @[LZD.scala 49:25]
  wire  _T_528; // @[LZD.scala 49:47]
  wire  _T_529; // @[LZD.scala 49:59]
  wire  _T_530; // @[LZD.scala 49:35]
  wire [2:0] _T_532; // @[Cat.scala 29:58]
  wire  _T_533; // @[Shift.scala 12:21]
  wire [2:0] _T_535; // @[LZD.scala 55:32]
  wire [2:0] _T_536; // @[LZD.scala 55:20]
  wire [3:0] _T_537; // @[Cat.scala 29:58]
  wire  _T_538; // @[Shift.scala 12:21]
  wire [3:0] _T_540; // @[LZD.scala 55:32]
  wire [3:0] _T_541; // @[LZD.scala 55:20]
  wire [4:0] _T_542; // @[Cat.scala 29:58]
  wire [4:0] _T_543; // @[convert.scala 21:22]
  wire [26:0] _T_544; // @[convert.scala 22:36]
  wire  _T_545; // @[Shift.scala 16:24]
  wire  _T_547; // @[Shift.scala 12:21]
  wire [10:0] _T_548; // @[Shift.scala 64:52]
  wire [26:0] _T_550; // @[Cat.scala 29:58]
  wire [26:0] _T_551; // @[Shift.scala 64:27]
  wire [3:0] _T_552; // @[Shift.scala 66:70]
  wire  _T_553; // @[Shift.scala 12:21]
  wire [18:0] _T_554; // @[Shift.scala 64:52]
  wire [26:0] _T_556; // @[Cat.scala 29:58]
  wire [26:0] _T_557; // @[Shift.scala 64:27]
  wire [2:0] _T_558; // @[Shift.scala 66:70]
  wire  _T_559; // @[Shift.scala 12:21]
  wire [22:0] _T_560; // @[Shift.scala 64:52]
  wire [26:0] _T_562; // @[Cat.scala 29:58]
  wire [26:0] _T_563; // @[Shift.scala 64:27]
  wire [1:0] _T_564; // @[Shift.scala 66:70]
  wire  _T_565; // @[Shift.scala 12:21]
  wire [24:0] _T_566; // @[Shift.scala 64:52]
  wire [26:0] _T_568; // @[Cat.scala 29:58]
  wire [26:0] _T_569; // @[Shift.scala 64:27]
  wire  _T_570; // @[Shift.scala 66:70]
  wire [25:0] _T_572; // @[Shift.scala 64:52]
  wire [26:0] _T_573; // @[Cat.scala 29:58]
  wire [26:0] _T_574; // @[Shift.scala 64:27]
  wire [26:0] _T_575; // @[Shift.scala 16:10]
  wire [2:0] _T_576; // @[convert.scala 23:34]
  wire [23:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_578; // @[convert.scala 25:26]
  wire [4:0] _T_580; // @[convert.scala 25:42]
  wire [2:0] _T_583; // @[convert.scala 26:67]
  wire [2:0] _T_584; // @[convert.scala 26:51]
  wire [8:0] _T_585; // @[Cat.scala 29:58]
  wire [28:0] _T_587; // @[convert.scala 29:56]
  wire  _T_588; // @[convert.scala 29:60]
  wire  _T_589; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_592; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [8:0] decB_scale; // @[convert.scala 32:24]
  wire  _T_601; // @[convert.scala 18:24]
  wire  _T_602; // @[convert.scala 18:40]
  wire  _T_603; // @[convert.scala 18:36]
  wire [27:0] _T_604; // @[convert.scala 19:24]
  wire [27:0] _T_605; // @[convert.scala 19:43]
  wire [27:0] _T_606; // @[convert.scala 19:39]
  wire [15:0] _T_607; // @[LZD.scala 43:32]
  wire [7:0] _T_608; // @[LZD.scala 43:32]
  wire [3:0] _T_609; // @[LZD.scala 43:32]
  wire [1:0] _T_610; // @[LZD.scala 43:32]
  wire  _T_611; // @[LZD.scala 39:14]
  wire  _T_612; // @[LZD.scala 39:21]
  wire  _T_613; // @[LZD.scala 39:30]
  wire  _T_614; // @[LZD.scala 39:27]
  wire  _T_615; // @[LZD.scala 39:25]
  wire [1:0] _T_616; // @[Cat.scala 29:58]
  wire [1:0] _T_617; // @[LZD.scala 44:32]
  wire  _T_618; // @[LZD.scala 39:14]
  wire  _T_619; // @[LZD.scala 39:21]
  wire  _T_620; // @[LZD.scala 39:30]
  wire  _T_621; // @[LZD.scala 39:27]
  wire  _T_622; // @[LZD.scala 39:25]
  wire [1:0] _T_623; // @[Cat.scala 29:58]
  wire  _T_624; // @[Shift.scala 12:21]
  wire  _T_625; // @[Shift.scala 12:21]
  wire  _T_626; // @[LZD.scala 49:16]
  wire  _T_627; // @[LZD.scala 49:27]
  wire  _T_628; // @[LZD.scala 49:25]
  wire  _T_629; // @[LZD.scala 49:47]
  wire  _T_630; // @[LZD.scala 49:59]
  wire  _T_631; // @[LZD.scala 49:35]
  wire [2:0] _T_633; // @[Cat.scala 29:58]
  wire [3:0] _T_634; // @[LZD.scala 44:32]
  wire [1:0] _T_635; // @[LZD.scala 43:32]
  wire  _T_636; // @[LZD.scala 39:14]
  wire  _T_637; // @[LZD.scala 39:21]
  wire  _T_638; // @[LZD.scala 39:30]
  wire  _T_639; // @[LZD.scala 39:27]
  wire  _T_640; // @[LZD.scala 39:25]
  wire [1:0] _T_641; // @[Cat.scala 29:58]
  wire [1:0] _T_642; // @[LZD.scala 44:32]
  wire  _T_643; // @[LZD.scala 39:14]
  wire  _T_644; // @[LZD.scala 39:21]
  wire  _T_645; // @[LZD.scala 39:30]
  wire  _T_646; // @[LZD.scala 39:27]
  wire  _T_647; // @[LZD.scala 39:25]
  wire [1:0] _T_648; // @[Cat.scala 29:58]
  wire  _T_649; // @[Shift.scala 12:21]
  wire  _T_650; // @[Shift.scala 12:21]
  wire  _T_651; // @[LZD.scala 49:16]
  wire  _T_652; // @[LZD.scala 49:27]
  wire  _T_653; // @[LZD.scala 49:25]
  wire  _T_654; // @[LZD.scala 49:47]
  wire  _T_655; // @[LZD.scala 49:59]
  wire  _T_656; // @[LZD.scala 49:35]
  wire [2:0] _T_658; // @[Cat.scala 29:58]
  wire  _T_659; // @[Shift.scala 12:21]
  wire  _T_660; // @[Shift.scala 12:21]
  wire  _T_661; // @[LZD.scala 49:16]
  wire  _T_662; // @[LZD.scala 49:27]
  wire  _T_663; // @[LZD.scala 49:25]
  wire [1:0] _T_664; // @[LZD.scala 49:47]
  wire [1:0] _T_665; // @[LZD.scala 49:59]
  wire [1:0] _T_666; // @[LZD.scala 49:35]
  wire [3:0] _T_668; // @[Cat.scala 29:58]
  wire [7:0] _T_669; // @[LZD.scala 44:32]
  wire [3:0] _T_670; // @[LZD.scala 43:32]
  wire [1:0] _T_671; // @[LZD.scala 43:32]
  wire  _T_672; // @[LZD.scala 39:14]
  wire  _T_673; // @[LZD.scala 39:21]
  wire  _T_674; // @[LZD.scala 39:30]
  wire  _T_675; // @[LZD.scala 39:27]
  wire  _T_676; // @[LZD.scala 39:25]
  wire [1:0] _T_677; // @[Cat.scala 29:58]
  wire [1:0] _T_678; // @[LZD.scala 44:32]
  wire  _T_679; // @[LZD.scala 39:14]
  wire  _T_680; // @[LZD.scala 39:21]
  wire  _T_681; // @[LZD.scala 39:30]
  wire  _T_682; // @[LZD.scala 39:27]
  wire  _T_683; // @[LZD.scala 39:25]
  wire [1:0] _T_684; // @[Cat.scala 29:58]
  wire  _T_685; // @[Shift.scala 12:21]
  wire  _T_686; // @[Shift.scala 12:21]
  wire  _T_687; // @[LZD.scala 49:16]
  wire  _T_688; // @[LZD.scala 49:27]
  wire  _T_689; // @[LZD.scala 49:25]
  wire  _T_690; // @[LZD.scala 49:47]
  wire  _T_691; // @[LZD.scala 49:59]
  wire  _T_692; // @[LZD.scala 49:35]
  wire [2:0] _T_694; // @[Cat.scala 29:58]
  wire [3:0] _T_695; // @[LZD.scala 44:32]
  wire [1:0] _T_696; // @[LZD.scala 43:32]
  wire  _T_697; // @[LZD.scala 39:14]
  wire  _T_698; // @[LZD.scala 39:21]
  wire  _T_699; // @[LZD.scala 39:30]
  wire  _T_700; // @[LZD.scala 39:27]
  wire  _T_701; // @[LZD.scala 39:25]
  wire [1:0] _T_702; // @[Cat.scala 29:58]
  wire [1:0] _T_703; // @[LZD.scala 44:32]
  wire  _T_704; // @[LZD.scala 39:14]
  wire  _T_705; // @[LZD.scala 39:21]
  wire  _T_706; // @[LZD.scala 39:30]
  wire  _T_707; // @[LZD.scala 39:27]
  wire  _T_708; // @[LZD.scala 39:25]
  wire [1:0] _T_709; // @[Cat.scala 29:58]
  wire  _T_710; // @[Shift.scala 12:21]
  wire  _T_711; // @[Shift.scala 12:21]
  wire  _T_712; // @[LZD.scala 49:16]
  wire  _T_713; // @[LZD.scala 49:27]
  wire  _T_714; // @[LZD.scala 49:25]
  wire  _T_715; // @[LZD.scala 49:47]
  wire  _T_716; // @[LZD.scala 49:59]
  wire  _T_717; // @[LZD.scala 49:35]
  wire [2:0] _T_719; // @[Cat.scala 29:58]
  wire  _T_720; // @[Shift.scala 12:21]
  wire  _T_721; // @[Shift.scala 12:21]
  wire  _T_722; // @[LZD.scala 49:16]
  wire  _T_723; // @[LZD.scala 49:27]
  wire  _T_724; // @[LZD.scala 49:25]
  wire [1:0] _T_725; // @[LZD.scala 49:47]
  wire [1:0] _T_726; // @[LZD.scala 49:59]
  wire [1:0] _T_727; // @[LZD.scala 49:35]
  wire [3:0] _T_729; // @[Cat.scala 29:58]
  wire  _T_730; // @[Shift.scala 12:21]
  wire  _T_731; // @[Shift.scala 12:21]
  wire  _T_732; // @[LZD.scala 49:16]
  wire  _T_733; // @[LZD.scala 49:27]
  wire  _T_734; // @[LZD.scala 49:25]
  wire [2:0] _T_735; // @[LZD.scala 49:47]
  wire [2:0] _T_736; // @[LZD.scala 49:59]
  wire [2:0] _T_737; // @[LZD.scala 49:35]
  wire [4:0] _T_739; // @[Cat.scala 29:58]
  wire [11:0] _T_740; // @[LZD.scala 44:32]
  wire [7:0] _T_741; // @[LZD.scala 43:32]
  wire [3:0] _T_742; // @[LZD.scala 43:32]
  wire [1:0] _T_743; // @[LZD.scala 43:32]
  wire  _T_744; // @[LZD.scala 39:14]
  wire  _T_745; // @[LZD.scala 39:21]
  wire  _T_746; // @[LZD.scala 39:30]
  wire  _T_747; // @[LZD.scala 39:27]
  wire  _T_748; // @[LZD.scala 39:25]
  wire [1:0] _T_749; // @[Cat.scala 29:58]
  wire [1:0] _T_750; // @[LZD.scala 44:32]
  wire  _T_751; // @[LZD.scala 39:14]
  wire  _T_752; // @[LZD.scala 39:21]
  wire  _T_753; // @[LZD.scala 39:30]
  wire  _T_754; // @[LZD.scala 39:27]
  wire  _T_755; // @[LZD.scala 39:25]
  wire [1:0] _T_756; // @[Cat.scala 29:58]
  wire  _T_757; // @[Shift.scala 12:21]
  wire  _T_758; // @[Shift.scala 12:21]
  wire  _T_759; // @[LZD.scala 49:16]
  wire  _T_760; // @[LZD.scala 49:27]
  wire  _T_761; // @[LZD.scala 49:25]
  wire  _T_762; // @[LZD.scala 49:47]
  wire  _T_763; // @[LZD.scala 49:59]
  wire  _T_764; // @[LZD.scala 49:35]
  wire [2:0] _T_766; // @[Cat.scala 29:58]
  wire [3:0] _T_767; // @[LZD.scala 44:32]
  wire [1:0] _T_768; // @[LZD.scala 43:32]
  wire  _T_769; // @[LZD.scala 39:14]
  wire  _T_770; // @[LZD.scala 39:21]
  wire  _T_771; // @[LZD.scala 39:30]
  wire  _T_772; // @[LZD.scala 39:27]
  wire  _T_773; // @[LZD.scala 39:25]
  wire [1:0] _T_774; // @[Cat.scala 29:58]
  wire [1:0] _T_775; // @[LZD.scala 44:32]
  wire  _T_776; // @[LZD.scala 39:14]
  wire  _T_777; // @[LZD.scala 39:21]
  wire  _T_778; // @[LZD.scala 39:30]
  wire  _T_779; // @[LZD.scala 39:27]
  wire  _T_780; // @[LZD.scala 39:25]
  wire [1:0] _T_781; // @[Cat.scala 29:58]
  wire  _T_782; // @[Shift.scala 12:21]
  wire  _T_783; // @[Shift.scala 12:21]
  wire  _T_784; // @[LZD.scala 49:16]
  wire  _T_785; // @[LZD.scala 49:27]
  wire  _T_786; // @[LZD.scala 49:25]
  wire  _T_787; // @[LZD.scala 49:47]
  wire  _T_788; // @[LZD.scala 49:59]
  wire  _T_789; // @[LZD.scala 49:35]
  wire [2:0] _T_791; // @[Cat.scala 29:58]
  wire  _T_792; // @[Shift.scala 12:21]
  wire  _T_793; // @[Shift.scala 12:21]
  wire  _T_794; // @[LZD.scala 49:16]
  wire  _T_795; // @[LZD.scala 49:27]
  wire  _T_796; // @[LZD.scala 49:25]
  wire [1:0] _T_797; // @[LZD.scala 49:47]
  wire [1:0] _T_798; // @[LZD.scala 49:59]
  wire [1:0] _T_799; // @[LZD.scala 49:35]
  wire [3:0] _T_801; // @[Cat.scala 29:58]
  wire [3:0] _T_802; // @[LZD.scala 44:32]
  wire [1:0] _T_803; // @[LZD.scala 43:32]
  wire  _T_804; // @[LZD.scala 39:14]
  wire  _T_805; // @[LZD.scala 39:21]
  wire  _T_806; // @[LZD.scala 39:30]
  wire  _T_807; // @[LZD.scala 39:27]
  wire  _T_808; // @[LZD.scala 39:25]
  wire [1:0] _T_809; // @[Cat.scala 29:58]
  wire [1:0] _T_810; // @[LZD.scala 44:32]
  wire  _T_811; // @[LZD.scala 39:14]
  wire  _T_812; // @[LZD.scala 39:21]
  wire  _T_813; // @[LZD.scala 39:30]
  wire  _T_814; // @[LZD.scala 39:27]
  wire  _T_815; // @[LZD.scala 39:25]
  wire [1:0] _T_816; // @[Cat.scala 29:58]
  wire  _T_817; // @[Shift.scala 12:21]
  wire  _T_818; // @[Shift.scala 12:21]
  wire  _T_819; // @[LZD.scala 49:16]
  wire  _T_820; // @[LZD.scala 49:27]
  wire  _T_821; // @[LZD.scala 49:25]
  wire  _T_822; // @[LZD.scala 49:47]
  wire  _T_823; // @[LZD.scala 49:59]
  wire  _T_824; // @[LZD.scala 49:35]
  wire [2:0] _T_826; // @[Cat.scala 29:58]
  wire  _T_827; // @[Shift.scala 12:21]
  wire [2:0] _T_829; // @[LZD.scala 55:32]
  wire [2:0] _T_830; // @[LZD.scala 55:20]
  wire [3:0] _T_831; // @[Cat.scala 29:58]
  wire  _T_832; // @[Shift.scala 12:21]
  wire [3:0] _T_834; // @[LZD.scala 55:32]
  wire [3:0] _T_835; // @[LZD.scala 55:20]
  wire [4:0] _T_836; // @[Cat.scala 29:58]
  wire [4:0] _T_837; // @[convert.scala 21:22]
  wire [26:0] _T_838; // @[convert.scala 22:36]
  wire  _T_839; // @[Shift.scala 16:24]
  wire  _T_841; // @[Shift.scala 12:21]
  wire [10:0] _T_842; // @[Shift.scala 64:52]
  wire [26:0] _T_844; // @[Cat.scala 29:58]
  wire [26:0] _T_845; // @[Shift.scala 64:27]
  wire [3:0] _T_846; // @[Shift.scala 66:70]
  wire  _T_847; // @[Shift.scala 12:21]
  wire [18:0] _T_848; // @[Shift.scala 64:52]
  wire [26:0] _T_850; // @[Cat.scala 29:58]
  wire [26:0] _T_851; // @[Shift.scala 64:27]
  wire [2:0] _T_852; // @[Shift.scala 66:70]
  wire  _T_853; // @[Shift.scala 12:21]
  wire [22:0] _T_854; // @[Shift.scala 64:52]
  wire [26:0] _T_856; // @[Cat.scala 29:58]
  wire [26:0] _T_857; // @[Shift.scala 64:27]
  wire [1:0] _T_858; // @[Shift.scala 66:70]
  wire  _T_859; // @[Shift.scala 12:21]
  wire [24:0] _T_860; // @[Shift.scala 64:52]
  wire [26:0] _T_862; // @[Cat.scala 29:58]
  wire [26:0] _T_863; // @[Shift.scala 64:27]
  wire  _T_864; // @[Shift.scala 66:70]
  wire [25:0] _T_866; // @[Shift.scala 64:52]
  wire [26:0] _T_867; // @[Cat.scala 29:58]
  wire [26:0] _T_868; // @[Shift.scala 64:27]
  wire [26:0] _T_869; // @[Shift.scala 16:10]
  wire [2:0] _T_870; // @[convert.scala 23:34]
  wire [23:0] decC_fraction; // @[convert.scala 24:34]
  wire  _T_872; // @[convert.scala 25:26]
  wire [4:0] _T_874; // @[convert.scala 25:42]
  wire [2:0] _T_877; // @[convert.scala 26:67]
  wire [2:0] _T_878; // @[convert.scala 26:51]
  wire [8:0] _T_879; // @[Cat.scala 29:58]
  wire [28:0] _T_881; // @[convert.scala 29:56]
  wire  _T_882; // @[convert.scala 29:60]
  wire  _T_883; // @[convert.scala 29:41]
  wire  decC_isNaR; // @[convert.scala 29:39]
  wire  _T_886; // @[convert.scala 30:19]
  wire  decC_isZero; // @[convert.scala 30:41]
  wire [8:0] decC_scale; // @[convert.scala 32:24]
  wire  _T_894; // @[PositFMA.scala 58:30]
  wire  outIsNaR; // @[PositFMA.scala 58:44]
  wire  _T_895; // @[PositFMA.scala 59:34]
  wire  _T_896; // @[PositFMA.scala 59:47]
  wire  _T_897; // @[PositFMA.scala 59:45]
  wire [25:0] _T_899; // @[Cat.scala 29:58]
  wire [25:0] sigA; // @[PositFMA.scala 59:76]
  wire  _T_900; // @[PositFMA.scala 60:34]
  wire  _T_901; // @[PositFMA.scala 60:47]
  wire  _T_902; // @[PositFMA.scala 60:45]
  wire [25:0] _T_904; // @[Cat.scala 29:58]
  wire [25:0] sigB; // @[PositFMA.scala 60:76]
  wire [51:0] _T_905; // @[PositFMA.scala 61:25]
  wire [51:0] sigP; // @[PositFMA.scala 61:33]
  wire [1:0] head2; // @[PositFMA.scala 62:28]
  wire  _T_906; // @[PositFMA.scala 63:31]
  wire  _T_907; // @[PositFMA.scala 63:25]
  wire  _T_908; // @[PositFMA.scala 63:42]
  wire  addTwo; // @[PositFMA.scala 63:35]
  wire  _T_909; // @[PositFMA.scala 65:23]
  wire  _T_910; // @[PositFMA.scala 65:49]
  wire  addOne; // @[PositFMA.scala 65:43]
  wire [1:0] _T_911; // @[Cat.scala 29:58]
  wire [2:0] expBias; // @[PositFMA.scala 66:39]
  wire  mulSign; // @[PositFMA.scala 67:28]
  wire [9:0] _T_912; // @[PositFMA.scala 69:30]
  wire [9:0] _GEN_12; // @[PositFMA.scala 69:44]
  wire [9:0] _T_914; // @[PositFMA.scala 69:44]
  wire [9:0] mulScale; // @[PositFMA.scala 69:44]
  wire [49:0] _T_915; // @[PositFMA.scala 72:29]
  wire [48:0] _T_916; // @[PositFMA.scala 73:29]
  wire [49:0] _T_917; // @[PositFMA.scala 73:48]
  wire [49:0] mulSigTmp; // @[PositFMA.scala 70:22]
  wire  _T_919; // @[PositFMA.scala 77:39]
  wire  _T_920; // @[PositFMA.scala 77:43]
  wire [48:0] _T_921; // @[PositFMA.scala 78:39]
  wire [50:0] mulSig; // @[Cat.scala 29:58]
  reg  outIsNaR_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg [50:0] mulSig_phase2; // @[Reg.scala 15:16]
  reg [63:0] _RAND_1;
  reg [23:0] addFrac_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [9:0] mulScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [8:0] addScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  addSign_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  addZero_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  inValid_phase2; // @[Valid.scala 117:22]
  reg [31:0] _RAND_7;
  wire  _T_947; // @[PositFMA.scala 107:29]
  wire  _T_948; // @[PositFMA.scala 107:47]
  wire  _T_949; // @[PositFMA.scala 107:45]
  wire [50:0] extAddSig; // @[Cat.scala 29:58]
  wire [9:0] _GEN_13; // @[PositFMA.scala 111:39]
  wire  mulGreater; // @[PositFMA.scala 111:39]
  wire [9:0] greaterScale; // @[PositFMA.scala 112:26]
  wire [9:0] smallerScale; // @[PositFMA.scala 113:26]
  wire [9:0] _T_953; // @[PositFMA.scala 114:36]
  wire [9:0] scaleDiff; // @[PositFMA.scala 114:36]
  wire [50:0] greaterSig; // @[PositFMA.scala 115:26]
  wire [50:0] smallerSigTmp; // @[PositFMA.scala 116:26]
  wire [9:0] _T_954; // @[PositFMA.scala 117:69]
  wire  _T_955; // @[Shift.scala 39:24]
  wire [5:0] _T_956; // @[Shift.scala 40:44]
  wire [18:0] _T_957; // @[Shift.scala 90:30]
  wire [31:0] _T_958; // @[Shift.scala 90:48]
  wire  _T_959; // @[Shift.scala 90:57]
  wire [18:0] _GEN_14; // @[Shift.scala 90:39]
  wire [18:0] _T_960; // @[Shift.scala 90:39]
  wire  _T_961; // @[Shift.scala 12:21]
  wire  _T_962; // @[Shift.scala 12:21]
  wire [31:0] _T_964; // @[Bitwise.scala 71:12]
  wire [50:0] _T_965; // @[Cat.scala 29:58]
  wire [50:0] _T_966; // @[Shift.scala 91:22]
  wire [4:0] _T_967; // @[Shift.scala 92:77]
  wire [34:0] _T_968; // @[Shift.scala 90:30]
  wire [15:0] _T_969; // @[Shift.scala 90:48]
  wire  _T_970; // @[Shift.scala 90:57]
  wire [34:0] _GEN_15; // @[Shift.scala 90:39]
  wire [34:0] _T_971; // @[Shift.scala 90:39]
  wire  _T_972; // @[Shift.scala 12:21]
  wire  _T_973; // @[Shift.scala 12:21]
  wire [15:0] _T_975; // @[Bitwise.scala 71:12]
  wire [50:0] _T_976; // @[Cat.scala 29:58]
  wire [50:0] _T_977; // @[Shift.scala 91:22]
  wire [3:0] _T_978; // @[Shift.scala 92:77]
  wire [42:0] _T_979; // @[Shift.scala 90:30]
  wire [7:0] _T_980; // @[Shift.scala 90:48]
  wire  _T_981; // @[Shift.scala 90:57]
  wire [42:0] _GEN_16; // @[Shift.scala 90:39]
  wire [42:0] _T_982; // @[Shift.scala 90:39]
  wire  _T_983; // @[Shift.scala 12:21]
  wire  _T_984; // @[Shift.scala 12:21]
  wire [7:0] _T_986; // @[Bitwise.scala 71:12]
  wire [50:0] _T_987; // @[Cat.scala 29:58]
  wire [50:0] _T_988; // @[Shift.scala 91:22]
  wire [2:0] _T_989; // @[Shift.scala 92:77]
  wire [46:0] _T_990; // @[Shift.scala 90:30]
  wire [3:0] _T_991; // @[Shift.scala 90:48]
  wire  _T_992; // @[Shift.scala 90:57]
  wire [46:0] _GEN_17; // @[Shift.scala 90:39]
  wire [46:0] _T_993; // @[Shift.scala 90:39]
  wire  _T_994; // @[Shift.scala 12:21]
  wire  _T_995; // @[Shift.scala 12:21]
  wire [3:0] _T_997; // @[Bitwise.scala 71:12]
  wire [50:0] _T_998; // @[Cat.scala 29:58]
  wire [50:0] _T_999; // @[Shift.scala 91:22]
  wire [1:0] _T_1000; // @[Shift.scala 92:77]
  wire [48:0] _T_1001; // @[Shift.scala 90:30]
  wire [1:0] _T_1002; // @[Shift.scala 90:48]
  wire  _T_1003; // @[Shift.scala 90:57]
  wire [48:0] _GEN_18; // @[Shift.scala 90:39]
  wire [48:0] _T_1004; // @[Shift.scala 90:39]
  wire  _T_1005; // @[Shift.scala 12:21]
  wire  _T_1006; // @[Shift.scala 12:21]
  wire [1:0] _T_1008; // @[Bitwise.scala 71:12]
  wire [50:0] _T_1009; // @[Cat.scala 29:58]
  wire [50:0] _T_1010; // @[Shift.scala 91:22]
  wire  _T_1011; // @[Shift.scala 92:77]
  wire [49:0] _T_1012; // @[Shift.scala 90:30]
  wire  _T_1013; // @[Shift.scala 90:48]
  wire [49:0] _GEN_19; // @[Shift.scala 90:39]
  wire [49:0] _T_1015; // @[Shift.scala 90:39]
  wire  _T_1017; // @[Shift.scala 12:21]
  wire [50:0] _T_1018; // @[Cat.scala 29:58]
  wire [50:0] _T_1019; // @[Shift.scala 91:22]
  wire [50:0] _T_1022; // @[Bitwise.scala 71:12]
  wire [50:0] smallerSig; // @[Shift.scala 39:10]
  wire [51:0] rawSumSig; // @[PositFMA.scala 118:34]
  wire  _T_1023; // @[PositFMA.scala 119:42]
  wire  _T_1024; // @[PositFMA.scala 119:46]
  wire  _T_1025; // @[PositFMA.scala 119:79]
  wire  sumSign; // @[PositFMA.scala 119:63]
  wire [50:0] _T_1027; // @[PositFMA.scala 120:50]
  wire [51:0] signSumSig; // @[Cat.scala 29:58]
  wire [50:0] _T_1028; // @[PositFMA.scala 124:33]
  wire [50:0] _T_1029; // @[PositFMA.scala 124:68]
  wire [50:0] sumXor; // @[PositFMA.scala 124:51]
  wire [31:0] _T_1030; // @[LZD.scala 43:32]
  wire [15:0] _T_1031; // @[LZD.scala 43:32]
  wire [7:0] _T_1032; // @[LZD.scala 43:32]
  wire [3:0] _T_1033; // @[LZD.scala 43:32]
  wire [1:0] _T_1034; // @[LZD.scala 43:32]
  wire  _T_1035; // @[LZD.scala 39:14]
  wire  _T_1036; // @[LZD.scala 39:21]
  wire  _T_1037; // @[LZD.scala 39:30]
  wire  _T_1038; // @[LZD.scala 39:27]
  wire  _T_1039; // @[LZD.scala 39:25]
  wire [1:0] _T_1040; // @[Cat.scala 29:58]
  wire [1:0] _T_1041; // @[LZD.scala 44:32]
  wire  _T_1042; // @[LZD.scala 39:14]
  wire  _T_1043; // @[LZD.scala 39:21]
  wire  _T_1044; // @[LZD.scala 39:30]
  wire  _T_1045; // @[LZD.scala 39:27]
  wire  _T_1046; // @[LZD.scala 39:25]
  wire [1:0] _T_1047; // @[Cat.scala 29:58]
  wire  _T_1048; // @[Shift.scala 12:21]
  wire  _T_1049; // @[Shift.scala 12:21]
  wire  _T_1050; // @[LZD.scala 49:16]
  wire  _T_1051; // @[LZD.scala 49:27]
  wire  _T_1052; // @[LZD.scala 49:25]
  wire  _T_1053; // @[LZD.scala 49:47]
  wire  _T_1054; // @[LZD.scala 49:59]
  wire  _T_1055; // @[LZD.scala 49:35]
  wire [2:0] _T_1057; // @[Cat.scala 29:58]
  wire [3:0] _T_1058; // @[LZD.scala 44:32]
  wire [1:0] _T_1059; // @[LZD.scala 43:32]
  wire  _T_1060; // @[LZD.scala 39:14]
  wire  _T_1061; // @[LZD.scala 39:21]
  wire  _T_1062; // @[LZD.scala 39:30]
  wire  _T_1063; // @[LZD.scala 39:27]
  wire  _T_1064; // @[LZD.scala 39:25]
  wire [1:0] _T_1065; // @[Cat.scala 29:58]
  wire [1:0] _T_1066; // @[LZD.scala 44:32]
  wire  _T_1067; // @[LZD.scala 39:14]
  wire  _T_1068; // @[LZD.scala 39:21]
  wire  _T_1069; // @[LZD.scala 39:30]
  wire  _T_1070; // @[LZD.scala 39:27]
  wire  _T_1071; // @[LZD.scala 39:25]
  wire [1:0] _T_1072; // @[Cat.scala 29:58]
  wire  _T_1073; // @[Shift.scala 12:21]
  wire  _T_1074; // @[Shift.scala 12:21]
  wire  _T_1075; // @[LZD.scala 49:16]
  wire  _T_1076; // @[LZD.scala 49:27]
  wire  _T_1077; // @[LZD.scala 49:25]
  wire  _T_1078; // @[LZD.scala 49:47]
  wire  _T_1079; // @[LZD.scala 49:59]
  wire  _T_1080; // @[LZD.scala 49:35]
  wire [2:0] _T_1082; // @[Cat.scala 29:58]
  wire  _T_1083; // @[Shift.scala 12:21]
  wire  _T_1084; // @[Shift.scala 12:21]
  wire  _T_1085; // @[LZD.scala 49:16]
  wire  _T_1086; // @[LZD.scala 49:27]
  wire  _T_1087; // @[LZD.scala 49:25]
  wire [1:0] _T_1088; // @[LZD.scala 49:47]
  wire [1:0] _T_1089; // @[LZD.scala 49:59]
  wire [1:0] _T_1090; // @[LZD.scala 49:35]
  wire [3:0] _T_1092; // @[Cat.scala 29:58]
  wire [7:0] _T_1093; // @[LZD.scala 44:32]
  wire [3:0] _T_1094; // @[LZD.scala 43:32]
  wire [1:0] _T_1095; // @[LZD.scala 43:32]
  wire  _T_1096; // @[LZD.scala 39:14]
  wire  _T_1097; // @[LZD.scala 39:21]
  wire  _T_1098; // @[LZD.scala 39:30]
  wire  _T_1099; // @[LZD.scala 39:27]
  wire  _T_1100; // @[LZD.scala 39:25]
  wire [1:0] _T_1101; // @[Cat.scala 29:58]
  wire [1:0] _T_1102; // @[LZD.scala 44:32]
  wire  _T_1103; // @[LZD.scala 39:14]
  wire  _T_1104; // @[LZD.scala 39:21]
  wire  _T_1105; // @[LZD.scala 39:30]
  wire  _T_1106; // @[LZD.scala 39:27]
  wire  _T_1107; // @[LZD.scala 39:25]
  wire [1:0] _T_1108; // @[Cat.scala 29:58]
  wire  _T_1109; // @[Shift.scala 12:21]
  wire  _T_1110; // @[Shift.scala 12:21]
  wire  _T_1111; // @[LZD.scala 49:16]
  wire  _T_1112; // @[LZD.scala 49:27]
  wire  _T_1113; // @[LZD.scala 49:25]
  wire  _T_1114; // @[LZD.scala 49:47]
  wire  _T_1115; // @[LZD.scala 49:59]
  wire  _T_1116; // @[LZD.scala 49:35]
  wire [2:0] _T_1118; // @[Cat.scala 29:58]
  wire [3:0] _T_1119; // @[LZD.scala 44:32]
  wire [1:0] _T_1120; // @[LZD.scala 43:32]
  wire  _T_1121; // @[LZD.scala 39:14]
  wire  _T_1122; // @[LZD.scala 39:21]
  wire  _T_1123; // @[LZD.scala 39:30]
  wire  _T_1124; // @[LZD.scala 39:27]
  wire  _T_1125; // @[LZD.scala 39:25]
  wire [1:0] _T_1126; // @[Cat.scala 29:58]
  wire [1:0] _T_1127; // @[LZD.scala 44:32]
  wire  _T_1128; // @[LZD.scala 39:14]
  wire  _T_1129; // @[LZD.scala 39:21]
  wire  _T_1130; // @[LZD.scala 39:30]
  wire  _T_1131; // @[LZD.scala 39:27]
  wire  _T_1132; // @[LZD.scala 39:25]
  wire [1:0] _T_1133; // @[Cat.scala 29:58]
  wire  _T_1134; // @[Shift.scala 12:21]
  wire  _T_1135; // @[Shift.scala 12:21]
  wire  _T_1136; // @[LZD.scala 49:16]
  wire  _T_1137; // @[LZD.scala 49:27]
  wire  _T_1138; // @[LZD.scala 49:25]
  wire  _T_1139; // @[LZD.scala 49:47]
  wire  _T_1140; // @[LZD.scala 49:59]
  wire  _T_1141; // @[LZD.scala 49:35]
  wire [2:0] _T_1143; // @[Cat.scala 29:58]
  wire  _T_1144; // @[Shift.scala 12:21]
  wire  _T_1145; // @[Shift.scala 12:21]
  wire  _T_1146; // @[LZD.scala 49:16]
  wire  _T_1147; // @[LZD.scala 49:27]
  wire  _T_1148; // @[LZD.scala 49:25]
  wire [1:0] _T_1149; // @[LZD.scala 49:47]
  wire [1:0] _T_1150; // @[LZD.scala 49:59]
  wire [1:0] _T_1151; // @[LZD.scala 49:35]
  wire [3:0] _T_1153; // @[Cat.scala 29:58]
  wire  _T_1154; // @[Shift.scala 12:21]
  wire  _T_1155; // @[Shift.scala 12:21]
  wire  _T_1156; // @[LZD.scala 49:16]
  wire  _T_1157; // @[LZD.scala 49:27]
  wire  _T_1158; // @[LZD.scala 49:25]
  wire [2:0] _T_1159; // @[LZD.scala 49:47]
  wire [2:0] _T_1160; // @[LZD.scala 49:59]
  wire [2:0] _T_1161; // @[LZD.scala 49:35]
  wire [4:0] _T_1163; // @[Cat.scala 29:58]
  wire [15:0] _T_1164; // @[LZD.scala 44:32]
  wire [7:0] _T_1165; // @[LZD.scala 43:32]
  wire [3:0] _T_1166; // @[LZD.scala 43:32]
  wire [1:0] _T_1167; // @[LZD.scala 43:32]
  wire  _T_1168; // @[LZD.scala 39:14]
  wire  _T_1169; // @[LZD.scala 39:21]
  wire  _T_1170; // @[LZD.scala 39:30]
  wire  _T_1171; // @[LZD.scala 39:27]
  wire  _T_1172; // @[LZD.scala 39:25]
  wire [1:0] _T_1173; // @[Cat.scala 29:58]
  wire [1:0] _T_1174; // @[LZD.scala 44:32]
  wire  _T_1175; // @[LZD.scala 39:14]
  wire  _T_1176; // @[LZD.scala 39:21]
  wire  _T_1177; // @[LZD.scala 39:30]
  wire  _T_1178; // @[LZD.scala 39:27]
  wire  _T_1179; // @[LZD.scala 39:25]
  wire [1:0] _T_1180; // @[Cat.scala 29:58]
  wire  _T_1181; // @[Shift.scala 12:21]
  wire  _T_1182; // @[Shift.scala 12:21]
  wire  _T_1183; // @[LZD.scala 49:16]
  wire  _T_1184; // @[LZD.scala 49:27]
  wire  _T_1185; // @[LZD.scala 49:25]
  wire  _T_1186; // @[LZD.scala 49:47]
  wire  _T_1187; // @[LZD.scala 49:59]
  wire  _T_1188; // @[LZD.scala 49:35]
  wire [2:0] _T_1190; // @[Cat.scala 29:58]
  wire [3:0] _T_1191; // @[LZD.scala 44:32]
  wire [1:0] _T_1192; // @[LZD.scala 43:32]
  wire  _T_1193; // @[LZD.scala 39:14]
  wire  _T_1194; // @[LZD.scala 39:21]
  wire  _T_1195; // @[LZD.scala 39:30]
  wire  _T_1196; // @[LZD.scala 39:27]
  wire  _T_1197; // @[LZD.scala 39:25]
  wire [1:0] _T_1198; // @[Cat.scala 29:58]
  wire [1:0] _T_1199; // @[LZD.scala 44:32]
  wire  _T_1200; // @[LZD.scala 39:14]
  wire  _T_1201; // @[LZD.scala 39:21]
  wire  _T_1202; // @[LZD.scala 39:30]
  wire  _T_1203; // @[LZD.scala 39:27]
  wire  _T_1204; // @[LZD.scala 39:25]
  wire [1:0] _T_1205; // @[Cat.scala 29:58]
  wire  _T_1206; // @[Shift.scala 12:21]
  wire  _T_1207; // @[Shift.scala 12:21]
  wire  _T_1208; // @[LZD.scala 49:16]
  wire  _T_1209; // @[LZD.scala 49:27]
  wire  _T_1210; // @[LZD.scala 49:25]
  wire  _T_1211; // @[LZD.scala 49:47]
  wire  _T_1212; // @[LZD.scala 49:59]
  wire  _T_1213; // @[LZD.scala 49:35]
  wire [2:0] _T_1215; // @[Cat.scala 29:58]
  wire  _T_1216; // @[Shift.scala 12:21]
  wire  _T_1217; // @[Shift.scala 12:21]
  wire  _T_1218; // @[LZD.scala 49:16]
  wire  _T_1219; // @[LZD.scala 49:27]
  wire  _T_1220; // @[LZD.scala 49:25]
  wire [1:0] _T_1221; // @[LZD.scala 49:47]
  wire [1:0] _T_1222; // @[LZD.scala 49:59]
  wire [1:0] _T_1223; // @[LZD.scala 49:35]
  wire [3:0] _T_1225; // @[Cat.scala 29:58]
  wire [7:0] _T_1226; // @[LZD.scala 44:32]
  wire [3:0] _T_1227; // @[LZD.scala 43:32]
  wire [1:0] _T_1228; // @[LZD.scala 43:32]
  wire  _T_1229; // @[LZD.scala 39:14]
  wire  _T_1230; // @[LZD.scala 39:21]
  wire  _T_1231; // @[LZD.scala 39:30]
  wire  _T_1232; // @[LZD.scala 39:27]
  wire  _T_1233; // @[LZD.scala 39:25]
  wire [1:0] _T_1234; // @[Cat.scala 29:58]
  wire [1:0] _T_1235; // @[LZD.scala 44:32]
  wire  _T_1236; // @[LZD.scala 39:14]
  wire  _T_1237; // @[LZD.scala 39:21]
  wire  _T_1238; // @[LZD.scala 39:30]
  wire  _T_1239; // @[LZD.scala 39:27]
  wire  _T_1240; // @[LZD.scala 39:25]
  wire [1:0] _T_1241; // @[Cat.scala 29:58]
  wire  _T_1242; // @[Shift.scala 12:21]
  wire  _T_1243; // @[Shift.scala 12:21]
  wire  _T_1244; // @[LZD.scala 49:16]
  wire  _T_1245; // @[LZD.scala 49:27]
  wire  _T_1246; // @[LZD.scala 49:25]
  wire  _T_1247; // @[LZD.scala 49:47]
  wire  _T_1248; // @[LZD.scala 49:59]
  wire  _T_1249; // @[LZD.scala 49:35]
  wire [2:0] _T_1251; // @[Cat.scala 29:58]
  wire [3:0] _T_1252; // @[LZD.scala 44:32]
  wire [1:0] _T_1253; // @[LZD.scala 43:32]
  wire  _T_1254; // @[LZD.scala 39:14]
  wire  _T_1255; // @[LZD.scala 39:21]
  wire  _T_1256; // @[LZD.scala 39:30]
  wire  _T_1257; // @[LZD.scala 39:27]
  wire  _T_1258; // @[LZD.scala 39:25]
  wire [1:0] _T_1259; // @[Cat.scala 29:58]
  wire [1:0] _T_1260; // @[LZD.scala 44:32]
  wire  _T_1261; // @[LZD.scala 39:14]
  wire  _T_1262; // @[LZD.scala 39:21]
  wire  _T_1263; // @[LZD.scala 39:30]
  wire  _T_1264; // @[LZD.scala 39:27]
  wire  _T_1265; // @[LZD.scala 39:25]
  wire [1:0] _T_1266; // @[Cat.scala 29:58]
  wire  _T_1267; // @[Shift.scala 12:21]
  wire  _T_1268; // @[Shift.scala 12:21]
  wire  _T_1269; // @[LZD.scala 49:16]
  wire  _T_1270; // @[LZD.scala 49:27]
  wire  _T_1271; // @[LZD.scala 49:25]
  wire  _T_1272; // @[LZD.scala 49:47]
  wire  _T_1273; // @[LZD.scala 49:59]
  wire  _T_1274; // @[LZD.scala 49:35]
  wire [2:0] _T_1276; // @[Cat.scala 29:58]
  wire  _T_1277; // @[Shift.scala 12:21]
  wire  _T_1278; // @[Shift.scala 12:21]
  wire  _T_1279; // @[LZD.scala 49:16]
  wire  _T_1280; // @[LZD.scala 49:27]
  wire  _T_1281; // @[LZD.scala 49:25]
  wire [1:0] _T_1282; // @[LZD.scala 49:47]
  wire [1:0] _T_1283; // @[LZD.scala 49:59]
  wire [1:0] _T_1284; // @[LZD.scala 49:35]
  wire [3:0] _T_1286; // @[Cat.scala 29:58]
  wire  _T_1287; // @[Shift.scala 12:21]
  wire  _T_1288; // @[Shift.scala 12:21]
  wire  _T_1289; // @[LZD.scala 49:16]
  wire  _T_1290; // @[LZD.scala 49:27]
  wire  _T_1291; // @[LZD.scala 49:25]
  wire [2:0] _T_1292; // @[LZD.scala 49:47]
  wire [2:0] _T_1293; // @[LZD.scala 49:59]
  wire [2:0] _T_1294; // @[LZD.scala 49:35]
  wire [4:0] _T_1296; // @[Cat.scala 29:58]
  wire  _T_1297; // @[Shift.scala 12:21]
  wire  _T_1298; // @[Shift.scala 12:21]
  wire  _T_1299; // @[LZD.scala 49:16]
  wire  _T_1300; // @[LZD.scala 49:27]
  wire  _T_1301; // @[LZD.scala 49:25]
  wire [3:0] _T_1302; // @[LZD.scala 49:47]
  wire [3:0] _T_1303; // @[LZD.scala 49:59]
  wire [3:0] _T_1304; // @[LZD.scala 49:35]
  wire [5:0] _T_1306; // @[Cat.scala 29:58]
  wire [18:0] _T_1307; // @[LZD.scala 44:32]
  wire [15:0] _T_1308; // @[LZD.scala 43:32]
  wire [7:0] _T_1309; // @[LZD.scala 43:32]
  wire [3:0] _T_1310; // @[LZD.scala 43:32]
  wire [1:0] _T_1311; // @[LZD.scala 43:32]
  wire  _T_1312; // @[LZD.scala 39:14]
  wire  _T_1313; // @[LZD.scala 39:21]
  wire  _T_1314; // @[LZD.scala 39:30]
  wire  _T_1315; // @[LZD.scala 39:27]
  wire  _T_1316; // @[LZD.scala 39:25]
  wire [1:0] _T_1317; // @[Cat.scala 29:58]
  wire [1:0] _T_1318; // @[LZD.scala 44:32]
  wire  _T_1319; // @[LZD.scala 39:14]
  wire  _T_1320; // @[LZD.scala 39:21]
  wire  _T_1321; // @[LZD.scala 39:30]
  wire  _T_1322; // @[LZD.scala 39:27]
  wire  _T_1323; // @[LZD.scala 39:25]
  wire [1:0] _T_1324; // @[Cat.scala 29:58]
  wire  _T_1325; // @[Shift.scala 12:21]
  wire  _T_1326; // @[Shift.scala 12:21]
  wire  _T_1327; // @[LZD.scala 49:16]
  wire  _T_1328; // @[LZD.scala 49:27]
  wire  _T_1329; // @[LZD.scala 49:25]
  wire  _T_1330; // @[LZD.scala 49:47]
  wire  _T_1331; // @[LZD.scala 49:59]
  wire  _T_1332; // @[LZD.scala 49:35]
  wire [2:0] _T_1334; // @[Cat.scala 29:58]
  wire [3:0] _T_1335; // @[LZD.scala 44:32]
  wire [1:0] _T_1336; // @[LZD.scala 43:32]
  wire  _T_1337; // @[LZD.scala 39:14]
  wire  _T_1338; // @[LZD.scala 39:21]
  wire  _T_1339; // @[LZD.scala 39:30]
  wire  _T_1340; // @[LZD.scala 39:27]
  wire  _T_1341; // @[LZD.scala 39:25]
  wire [1:0] _T_1342; // @[Cat.scala 29:58]
  wire [1:0] _T_1343; // @[LZD.scala 44:32]
  wire  _T_1344; // @[LZD.scala 39:14]
  wire  _T_1345; // @[LZD.scala 39:21]
  wire  _T_1346; // @[LZD.scala 39:30]
  wire  _T_1347; // @[LZD.scala 39:27]
  wire  _T_1348; // @[LZD.scala 39:25]
  wire [1:0] _T_1349; // @[Cat.scala 29:58]
  wire  _T_1350; // @[Shift.scala 12:21]
  wire  _T_1351; // @[Shift.scala 12:21]
  wire  _T_1352; // @[LZD.scala 49:16]
  wire  _T_1353; // @[LZD.scala 49:27]
  wire  _T_1354; // @[LZD.scala 49:25]
  wire  _T_1355; // @[LZD.scala 49:47]
  wire  _T_1356; // @[LZD.scala 49:59]
  wire  _T_1357; // @[LZD.scala 49:35]
  wire [2:0] _T_1359; // @[Cat.scala 29:58]
  wire  _T_1360; // @[Shift.scala 12:21]
  wire  _T_1361; // @[Shift.scala 12:21]
  wire  _T_1362; // @[LZD.scala 49:16]
  wire  _T_1363; // @[LZD.scala 49:27]
  wire  _T_1364; // @[LZD.scala 49:25]
  wire [1:0] _T_1365; // @[LZD.scala 49:47]
  wire [1:0] _T_1366; // @[LZD.scala 49:59]
  wire [1:0] _T_1367; // @[LZD.scala 49:35]
  wire [3:0] _T_1369; // @[Cat.scala 29:58]
  wire [7:0] _T_1370; // @[LZD.scala 44:32]
  wire [3:0] _T_1371; // @[LZD.scala 43:32]
  wire [1:0] _T_1372; // @[LZD.scala 43:32]
  wire  _T_1373; // @[LZD.scala 39:14]
  wire  _T_1374; // @[LZD.scala 39:21]
  wire  _T_1375; // @[LZD.scala 39:30]
  wire  _T_1376; // @[LZD.scala 39:27]
  wire  _T_1377; // @[LZD.scala 39:25]
  wire [1:0] _T_1378; // @[Cat.scala 29:58]
  wire [1:0] _T_1379; // @[LZD.scala 44:32]
  wire  _T_1380; // @[LZD.scala 39:14]
  wire  _T_1381; // @[LZD.scala 39:21]
  wire  _T_1382; // @[LZD.scala 39:30]
  wire  _T_1383; // @[LZD.scala 39:27]
  wire  _T_1384; // @[LZD.scala 39:25]
  wire [1:0] _T_1385; // @[Cat.scala 29:58]
  wire  _T_1386; // @[Shift.scala 12:21]
  wire  _T_1387; // @[Shift.scala 12:21]
  wire  _T_1388; // @[LZD.scala 49:16]
  wire  _T_1389; // @[LZD.scala 49:27]
  wire  _T_1390; // @[LZD.scala 49:25]
  wire  _T_1391; // @[LZD.scala 49:47]
  wire  _T_1392; // @[LZD.scala 49:59]
  wire  _T_1393; // @[LZD.scala 49:35]
  wire [2:0] _T_1395; // @[Cat.scala 29:58]
  wire [3:0] _T_1396; // @[LZD.scala 44:32]
  wire [1:0] _T_1397; // @[LZD.scala 43:32]
  wire  _T_1398; // @[LZD.scala 39:14]
  wire  _T_1399; // @[LZD.scala 39:21]
  wire  _T_1400; // @[LZD.scala 39:30]
  wire  _T_1401; // @[LZD.scala 39:27]
  wire  _T_1402; // @[LZD.scala 39:25]
  wire [1:0] _T_1403; // @[Cat.scala 29:58]
  wire [1:0] _T_1404; // @[LZD.scala 44:32]
  wire  _T_1405; // @[LZD.scala 39:14]
  wire  _T_1406; // @[LZD.scala 39:21]
  wire  _T_1407; // @[LZD.scala 39:30]
  wire  _T_1408; // @[LZD.scala 39:27]
  wire  _T_1409; // @[LZD.scala 39:25]
  wire [1:0] _T_1410; // @[Cat.scala 29:58]
  wire  _T_1411; // @[Shift.scala 12:21]
  wire  _T_1412; // @[Shift.scala 12:21]
  wire  _T_1413; // @[LZD.scala 49:16]
  wire  _T_1414; // @[LZD.scala 49:27]
  wire  _T_1415; // @[LZD.scala 49:25]
  wire  _T_1416; // @[LZD.scala 49:47]
  wire  _T_1417; // @[LZD.scala 49:59]
  wire  _T_1418; // @[LZD.scala 49:35]
  wire [2:0] _T_1420; // @[Cat.scala 29:58]
  wire  _T_1421; // @[Shift.scala 12:21]
  wire  _T_1422; // @[Shift.scala 12:21]
  wire  _T_1423; // @[LZD.scala 49:16]
  wire  _T_1424; // @[LZD.scala 49:27]
  wire  _T_1425; // @[LZD.scala 49:25]
  wire [1:0] _T_1426; // @[LZD.scala 49:47]
  wire [1:0] _T_1427; // @[LZD.scala 49:59]
  wire [1:0] _T_1428; // @[LZD.scala 49:35]
  wire [3:0] _T_1430; // @[Cat.scala 29:58]
  wire  _T_1431; // @[Shift.scala 12:21]
  wire  _T_1432; // @[Shift.scala 12:21]
  wire  _T_1433; // @[LZD.scala 49:16]
  wire  _T_1434; // @[LZD.scala 49:27]
  wire  _T_1435; // @[LZD.scala 49:25]
  wire [2:0] _T_1436; // @[LZD.scala 49:47]
  wire [2:0] _T_1437; // @[LZD.scala 49:59]
  wire [2:0] _T_1438; // @[LZD.scala 49:35]
  wire [4:0] _T_1440; // @[Cat.scala 29:58]
  wire [2:0] _T_1441; // @[LZD.scala 44:32]
  wire [1:0] _T_1442; // @[LZD.scala 43:32]
  wire  _T_1443; // @[LZD.scala 39:14]
  wire  _T_1444; // @[LZD.scala 39:21]
  wire  _T_1445; // @[LZD.scala 39:30]
  wire  _T_1446; // @[LZD.scala 39:27]
  wire  _T_1447; // @[LZD.scala 39:25]
  wire [1:0] _T_1448; // @[Cat.scala 29:58]
  wire  _T_1449; // @[LZD.scala 44:32]
  wire  _T_1451; // @[Shift.scala 12:21]
  wire  _T_1453; // @[LZD.scala 55:32]
  wire  _T_1454; // @[LZD.scala 55:20]
  wire  _T_1456; // @[Shift.scala 12:21]
  wire [3:0] _T_1459; // @[Cat.scala 29:58]
  wire [3:0] _T_1460; // @[LZD.scala 55:32]
  wire [3:0] _T_1461; // @[LZD.scala 55:20]
  wire [4:0] _T_1462; // @[Cat.scala 29:58]
  wire  _T_1463; // @[Shift.scala 12:21]
  wire [4:0] _T_1465; // @[LZD.scala 55:32]
  wire [4:0] _T_1466; // @[LZD.scala 55:20]
  wire [5:0] sumLZD; // @[Cat.scala 29:58]
  wire [5:0] shiftValue; // @[PositFMA.scala 126:24]
  wire [49:0] _T_1467; // @[PositFMA.scala 127:38]
  wire  _T_1468; // @[Shift.scala 16:24]
  wire  _T_1470; // @[Shift.scala 12:21]
  wire [17:0] _T_1471; // @[Shift.scala 64:52]
  wire [49:0] _T_1473; // @[Cat.scala 29:58]
  wire [49:0] _T_1474; // @[Shift.scala 64:27]
  wire [4:0] _T_1475; // @[Shift.scala 66:70]
  wire  _T_1476; // @[Shift.scala 12:21]
  wire [33:0] _T_1477; // @[Shift.scala 64:52]
  wire [49:0] _T_1479; // @[Cat.scala 29:58]
  wire [49:0] _T_1480; // @[Shift.scala 64:27]
  wire [3:0] _T_1481; // @[Shift.scala 66:70]
  wire  _T_1482; // @[Shift.scala 12:21]
  wire [41:0] _T_1483; // @[Shift.scala 64:52]
  wire [49:0] _T_1485; // @[Cat.scala 29:58]
  wire [49:0] _T_1486; // @[Shift.scala 64:27]
  wire [2:0] _T_1487; // @[Shift.scala 66:70]
  wire  _T_1488; // @[Shift.scala 12:21]
  wire [45:0] _T_1489; // @[Shift.scala 64:52]
  wire [49:0] _T_1491; // @[Cat.scala 29:58]
  wire [49:0] _T_1492; // @[Shift.scala 64:27]
  wire [1:0] _T_1493; // @[Shift.scala 66:70]
  wire  _T_1494; // @[Shift.scala 12:21]
  wire [47:0] _T_1495; // @[Shift.scala 64:52]
  wire [49:0] _T_1497; // @[Cat.scala 29:58]
  wire [49:0] _T_1498; // @[Shift.scala 64:27]
  wire  _T_1499; // @[Shift.scala 66:70]
  wire [48:0] _T_1501; // @[Shift.scala 64:52]
  wire [49:0] _T_1502; // @[Cat.scala 29:58]
  wire [49:0] _T_1503; // @[Shift.scala 64:27]
  wire [49:0] normalFracTmp; // @[Shift.scala 16:10]
  wire [9:0] _T_1505; // @[PositFMA.scala 130:36]
  wire [9:0] _T_1506; // @[PositFMA.scala 130:36]
  wire [6:0] _T_1507; // @[Cat.scala 29:58]
  wire [6:0] _T_1508; // @[PositFMA.scala 130:61]
  wire [9:0] _GEN_20; // @[PositFMA.scala 130:42]
  wire [9:0] _T_1510; // @[PositFMA.scala 130:42]
  wire [9:0] sumScale; // @[PositFMA.scala 130:42]
  wire [23:0] sumFrac; // @[PositFMA.scala 131:41]
  wire [25:0] grsTmp; // @[PositFMA.scala 134:41]
  wire [1:0] _T_1511; // @[PositFMA.scala 137:40]
  wire [23:0] _T_1512; // @[PositFMA.scala 137:56]
  wire  _T_1513; // @[PositFMA.scala 137:60]
  wire  underflow; // @[PositFMA.scala 144:32]
  wire  overflow; // @[PositFMA.scala 145:32]
  wire  _T_1514; // @[PositFMA.scala 154:32]
  wire  decF_isZero; // @[PositFMA.scala 154:20]
  wire [9:0] _T_1516; // @[Mux.scala 87:16]
  wire [9:0] _T_1517; // @[Mux.scala 87:16]
  wire [8:0] _GEN_21; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  wire [8:0] decF_scale; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  wire [2:0] _T_1518; // @[convert.scala 46:61]
  wire [2:0] _T_1519; // @[convert.scala 46:52]
  wire [2:0] _T_1521; // @[convert.scala 46:42]
  wire [5:0] _T_1522; // @[convert.scala 48:34]
  wire  _T_1523; // @[convert.scala 49:36]
  wire [5:0] _T_1525; // @[convert.scala 50:36]
  wire [5:0] _T_1526; // @[convert.scala 50:36]
  wire [5:0] _T_1527; // @[convert.scala 50:28]
  wire  _T_1528; // @[convert.scala 51:31]
  wire  _T_1529; // @[convert.scala 52:43]
  wire [31:0] _T_1533; // @[Cat.scala 29:58]
  wire [5:0] _T_1534; // @[Shift.scala 39:17]
  wire  _T_1535; // @[Shift.scala 39:24]
  wire [4:0] _T_1536; // @[Shift.scala 40:44]
  wire [15:0] _T_1537; // @[Shift.scala 90:30]
  wire [15:0] _T_1538; // @[Shift.scala 90:48]
  wire  _T_1539; // @[Shift.scala 90:57]
  wire [15:0] _GEN_22; // @[Shift.scala 90:39]
  wire [15:0] _T_1540; // @[Shift.scala 90:39]
  wire  _T_1541; // @[Shift.scala 12:21]
  wire  _T_1542; // @[Shift.scala 12:21]
  wire [15:0] _T_1544; // @[Bitwise.scala 71:12]
  wire [31:0] _T_1545; // @[Cat.scala 29:58]
  wire [31:0] _T_1546; // @[Shift.scala 91:22]
  wire [3:0] _T_1547; // @[Shift.scala 92:77]
  wire [23:0] _T_1548; // @[Shift.scala 90:30]
  wire [7:0] _T_1549; // @[Shift.scala 90:48]
  wire  _T_1550; // @[Shift.scala 90:57]
  wire [23:0] _GEN_23; // @[Shift.scala 90:39]
  wire [23:0] _T_1551; // @[Shift.scala 90:39]
  wire  _T_1552; // @[Shift.scala 12:21]
  wire  _T_1553; // @[Shift.scala 12:21]
  wire [7:0] _T_1555; // @[Bitwise.scala 71:12]
  wire [31:0] _T_1556; // @[Cat.scala 29:58]
  wire [31:0] _T_1557; // @[Shift.scala 91:22]
  wire [2:0] _T_1558; // @[Shift.scala 92:77]
  wire [27:0] _T_1559; // @[Shift.scala 90:30]
  wire [3:0] _T_1560; // @[Shift.scala 90:48]
  wire  _T_1561; // @[Shift.scala 90:57]
  wire [27:0] _GEN_24; // @[Shift.scala 90:39]
  wire [27:0] _T_1562; // @[Shift.scala 90:39]
  wire  _T_1563; // @[Shift.scala 12:21]
  wire  _T_1564; // @[Shift.scala 12:21]
  wire [3:0] _T_1566; // @[Bitwise.scala 71:12]
  wire [31:0] _T_1567; // @[Cat.scala 29:58]
  wire [31:0] _T_1568; // @[Shift.scala 91:22]
  wire [1:0] _T_1569; // @[Shift.scala 92:77]
  wire [29:0] _T_1570; // @[Shift.scala 90:30]
  wire [1:0] _T_1571; // @[Shift.scala 90:48]
  wire  _T_1572; // @[Shift.scala 90:57]
  wire [29:0] _GEN_25; // @[Shift.scala 90:39]
  wire [29:0] _T_1573; // @[Shift.scala 90:39]
  wire  _T_1574; // @[Shift.scala 12:21]
  wire  _T_1575; // @[Shift.scala 12:21]
  wire [1:0] _T_1577; // @[Bitwise.scala 71:12]
  wire [31:0] _T_1578; // @[Cat.scala 29:58]
  wire [31:0] _T_1579; // @[Shift.scala 91:22]
  wire  _T_1580; // @[Shift.scala 92:77]
  wire [30:0] _T_1581; // @[Shift.scala 90:30]
  wire  _T_1582; // @[Shift.scala 90:48]
  wire [30:0] _GEN_26; // @[Shift.scala 90:39]
  wire [30:0] _T_1584; // @[Shift.scala 90:39]
  wire  _T_1586; // @[Shift.scala 12:21]
  wire [31:0] _T_1587; // @[Cat.scala 29:58]
  wire [31:0] _T_1588; // @[Shift.scala 91:22]
  wire [31:0] _T_1591; // @[Bitwise.scala 71:12]
  wire [31:0] _T_1592; // @[Shift.scala 39:10]
  wire  _T_1593; // @[convert.scala 55:31]
  wire  _T_1594; // @[convert.scala 56:31]
  wire  _T_1595; // @[convert.scala 57:31]
  wire  _T_1596; // @[convert.scala 58:31]
  wire [28:0] _T_1597; // @[convert.scala 59:69]
  wire  _T_1598; // @[convert.scala 59:81]
  wire  _T_1599; // @[convert.scala 59:50]
  wire  _T_1601; // @[convert.scala 60:81]
  wire  _T_1602; // @[convert.scala 61:44]
  wire  _T_1603; // @[convert.scala 61:52]
  wire  _T_1604; // @[convert.scala 61:36]
  wire  _T_1605; // @[convert.scala 62:63]
  wire  _T_1606; // @[convert.scala 62:103]
  wire  _T_1607; // @[convert.scala 62:60]
  wire [28:0] _GEN_27; // @[convert.scala 63:56]
  wire [28:0] _T_1610; // @[convert.scala 63:56]
  wire [29:0] _T_1611; // @[Cat.scala 29:58]
  reg  _T_1615; // @[Valid.scala 117:22]
  reg [31:0] _RAND_8;
  reg [29:0] _T_1619; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  assign _T = io_fmaOp[1]; // @[PositFMA.scala 47:36]
  assign _T_2 = _T ? 30'h3fffffff : 30'h0; // @[Bitwise.scala 71:12]
  assign _T_3 = _T_2 ^ io_A; // @[PositFMA.scala 47:41]
  assign _GEN_10 = {{29'd0}, _T}; // @[PositFMA.scala 47:49]
  assign realA = _T_3 + _GEN_10; // @[PositFMA.scala 47:49]
  assign _T_6 = io_fmaOp[0]; // @[PositFMA.scala 48:36]
  assign _T_8 = _T_6 ? 30'h3fffffff : 30'h0; // @[Bitwise.scala 71:12]
  assign _T_9 = _T_8 ^ io_C; // @[PositFMA.scala 48:41]
  assign _GEN_11 = {{29'd0}, _T_6}; // @[PositFMA.scala 48:49]
  assign realC = _T_9 + _GEN_11; // @[PositFMA.scala 48:49]
  assign _T_13 = realA[29]; // @[convert.scala 18:24]
  assign _T_14 = realA[28]; // @[convert.scala 18:40]
  assign _T_15 = _T_13 ^ _T_14; // @[convert.scala 18:36]
  assign _T_16 = realA[28:1]; // @[convert.scala 19:24]
  assign _T_17 = realA[27:0]; // @[convert.scala 19:43]
  assign _T_18 = _T_16 ^ _T_17; // @[convert.scala 19:39]
  assign _T_19 = _T_18[27:12]; // @[LZD.scala 43:32]
  assign _T_20 = _T_19[15:8]; // @[LZD.scala 43:32]
  assign _T_21 = _T_20[7:4]; // @[LZD.scala 43:32]
  assign _T_22 = _T_21[3:2]; // @[LZD.scala 43:32]
  assign _T_23 = _T_22 != 2'h0; // @[LZD.scala 39:14]
  assign _T_24 = _T_22[1]; // @[LZD.scala 39:21]
  assign _T_25 = _T_22[0]; // @[LZD.scala 39:30]
  assign _T_26 = ~ _T_25; // @[LZD.scala 39:27]
  assign _T_27 = _T_24 | _T_26; // @[LZD.scala 39:25]
  assign _T_28 = {_T_23,_T_27}; // @[Cat.scala 29:58]
  assign _T_29 = _T_21[1:0]; // @[LZD.scala 44:32]
  assign _T_30 = _T_29 != 2'h0; // @[LZD.scala 39:14]
  assign _T_31 = _T_29[1]; // @[LZD.scala 39:21]
  assign _T_32 = _T_29[0]; // @[LZD.scala 39:30]
  assign _T_33 = ~ _T_32; // @[LZD.scala 39:27]
  assign _T_34 = _T_31 | _T_33; // @[LZD.scala 39:25]
  assign _T_35 = {_T_30,_T_34}; // @[Cat.scala 29:58]
  assign _T_36 = _T_28[1]; // @[Shift.scala 12:21]
  assign _T_37 = _T_35[1]; // @[Shift.scala 12:21]
  assign _T_38 = _T_36 | _T_37; // @[LZD.scala 49:16]
  assign _T_39 = ~ _T_37; // @[LZD.scala 49:27]
  assign _T_40 = _T_36 | _T_39; // @[LZD.scala 49:25]
  assign _T_41 = _T_28[0:0]; // @[LZD.scala 49:47]
  assign _T_42 = _T_35[0:0]; // @[LZD.scala 49:59]
  assign _T_43 = _T_36 ? _T_41 : _T_42; // @[LZD.scala 49:35]
  assign _T_45 = {_T_38,_T_40,_T_43}; // @[Cat.scala 29:58]
  assign _T_46 = _T_20[3:0]; // @[LZD.scala 44:32]
  assign _T_47 = _T_46[3:2]; // @[LZD.scala 43:32]
  assign _T_48 = _T_47 != 2'h0; // @[LZD.scala 39:14]
  assign _T_49 = _T_47[1]; // @[LZD.scala 39:21]
  assign _T_50 = _T_47[0]; // @[LZD.scala 39:30]
  assign _T_51 = ~ _T_50; // @[LZD.scala 39:27]
  assign _T_52 = _T_49 | _T_51; // @[LZD.scala 39:25]
  assign _T_53 = {_T_48,_T_52}; // @[Cat.scala 29:58]
  assign _T_54 = _T_46[1:0]; // @[LZD.scala 44:32]
  assign _T_55 = _T_54 != 2'h0; // @[LZD.scala 39:14]
  assign _T_56 = _T_54[1]; // @[LZD.scala 39:21]
  assign _T_57 = _T_54[0]; // @[LZD.scala 39:30]
  assign _T_58 = ~ _T_57; // @[LZD.scala 39:27]
  assign _T_59 = _T_56 | _T_58; // @[LZD.scala 39:25]
  assign _T_60 = {_T_55,_T_59}; // @[Cat.scala 29:58]
  assign _T_61 = _T_53[1]; // @[Shift.scala 12:21]
  assign _T_62 = _T_60[1]; // @[Shift.scala 12:21]
  assign _T_63 = _T_61 | _T_62; // @[LZD.scala 49:16]
  assign _T_64 = ~ _T_62; // @[LZD.scala 49:27]
  assign _T_65 = _T_61 | _T_64; // @[LZD.scala 49:25]
  assign _T_66 = _T_53[0:0]; // @[LZD.scala 49:47]
  assign _T_67 = _T_60[0:0]; // @[LZD.scala 49:59]
  assign _T_68 = _T_61 ? _T_66 : _T_67; // @[LZD.scala 49:35]
  assign _T_70 = {_T_63,_T_65,_T_68}; // @[Cat.scala 29:58]
  assign _T_71 = _T_45[2]; // @[Shift.scala 12:21]
  assign _T_72 = _T_70[2]; // @[Shift.scala 12:21]
  assign _T_73 = _T_71 | _T_72; // @[LZD.scala 49:16]
  assign _T_74 = ~ _T_72; // @[LZD.scala 49:27]
  assign _T_75 = _T_71 | _T_74; // @[LZD.scala 49:25]
  assign _T_76 = _T_45[1:0]; // @[LZD.scala 49:47]
  assign _T_77 = _T_70[1:0]; // @[LZD.scala 49:59]
  assign _T_78 = _T_71 ? _T_76 : _T_77; // @[LZD.scala 49:35]
  assign _T_80 = {_T_73,_T_75,_T_78}; // @[Cat.scala 29:58]
  assign _T_81 = _T_19[7:0]; // @[LZD.scala 44:32]
  assign _T_82 = _T_81[7:4]; // @[LZD.scala 43:32]
  assign _T_83 = _T_82[3:2]; // @[LZD.scala 43:32]
  assign _T_84 = _T_83 != 2'h0; // @[LZD.scala 39:14]
  assign _T_85 = _T_83[1]; // @[LZD.scala 39:21]
  assign _T_86 = _T_83[0]; // @[LZD.scala 39:30]
  assign _T_87 = ~ _T_86; // @[LZD.scala 39:27]
  assign _T_88 = _T_85 | _T_87; // @[LZD.scala 39:25]
  assign _T_89 = {_T_84,_T_88}; // @[Cat.scala 29:58]
  assign _T_90 = _T_82[1:0]; // @[LZD.scala 44:32]
  assign _T_91 = _T_90 != 2'h0; // @[LZD.scala 39:14]
  assign _T_92 = _T_90[1]; // @[LZD.scala 39:21]
  assign _T_93 = _T_90[0]; // @[LZD.scala 39:30]
  assign _T_94 = ~ _T_93; // @[LZD.scala 39:27]
  assign _T_95 = _T_92 | _T_94; // @[LZD.scala 39:25]
  assign _T_96 = {_T_91,_T_95}; // @[Cat.scala 29:58]
  assign _T_97 = _T_89[1]; // @[Shift.scala 12:21]
  assign _T_98 = _T_96[1]; // @[Shift.scala 12:21]
  assign _T_99 = _T_97 | _T_98; // @[LZD.scala 49:16]
  assign _T_100 = ~ _T_98; // @[LZD.scala 49:27]
  assign _T_101 = _T_97 | _T_100; // @[LZD.scala 49:25]
  assign _T_102 = _T_89[0:0]; // @[LZD.scala 49:47]
  assign _T_103 = _T_96[0:0]; // @[LZD.scala 49:59]
  assign _T_104 = _T_97 ? _T_102 : _T_103; // @[LZD.scala 49:35]
  assign _T_106 = {_T_99,_T_101,_T_104}; // @[Cat.scala 29:58]
  assign _T_107 = _T_81[3:0]; // @[LZD.scala 44:32]
  assign _T_108 = _T_107[3:2]; // @[LZD.scala 43:32]
  assign _T_109 = _T_108 != 2'h0; // @[LZD.scala 39:14]
  assign _T_110 = _T_108[1]; // @[LZD.scala 39:21]
  assign _T_111 = _T_108[0]; // @[LZD.scala 39:30]
  assign _T_112 = ~ _T_111; // @[LZD.scala 39:27]
  assign _T_113 = _T_110 | _T_112; // @[LZD.scala 39:25]
  assign _T_114 = {_T_109,_T_113}; // @[Cat.scala 29:58]
  assign _T_115 = _T_107[1:0]; // @[LZD.scala 44:32]
  assign _T_116 = _T_115 != 2'h0; // @[LZD.scala 39:14]
  assign _T_117 = _T_115[1]; // @[LZD.scala 39:21]
  assign _T_118 = _T_115[0]; // @[LZD.scala 39:30]
  assign _T_119 = ~ _T_118; // @[LZD.scala 39:27]
  assign _T_120 = _T_117 | _T_119; // @[LZD.scala 39:25]
  assign _T_121 = {_T_116,_T_120}; // @[Cat.scala 29:58]
  assign _T_122 = _T_114[1]; // @[Shift.scala 12:21]
  assign _T_123 = _T_121[1]; // @[Shift.scala 12:21]
  assign _T_124 = _T_122 | _T_123; // @[LZD.scala 49:16]
  assign _T_125 = ~ _T_123; // @[LZD.scala 49:27]
  assign _T_126 = _T_122 | _T_125; // @[LZD.scala 49:25]
  assign _T_127 = _T_114[0:0]; // @[LZD.scala 49:47]
  assign _T_128 = _T_121[0:0]; // @[LZD.scala 49:59]
  assign _T_129 = _T_122 ? _T_127 : _T_128; // @[LZD.scala 49:35]
  assign _T_131 = {_T_124,_T_126,_T_129}; // @[Cat.scala 29:58]
  assign _T_132 = _T_106[2]; // @[Shift.scala 12:21]
  assign _T_133 = _T_131[2]; // @[Shift.scala 12:21]
  assign _T_134 = _T_132 | _T_133; // @[LZD.scala 49:16]
  assign _T_135 = ~ _T_133; // @[LZD.scala 49:27]
  assign _T_136 = _T_132 | _T_135; // @[LZD.scala 49:25]
  assign _T_137 = _T_106[1:0]; // @[LZD.scala 49:47]
  assign _T_138 = _T_131[1:0]; // @[LZD.scala 49:59]
  assign _T_139 = _T_132 ? _T_137 : _T_138; // @[LZD.scala 49:35]
  assign _T_141 = {_T_134,_T_136,_T_139}; // @[Cat.scala 29:58]
  assign _T_142 = _T_80[3]; // @[Shift.scala 12:21]
  assign _T_143 = _T_141[3]; // @[Shift.scala 12:21]
  assign _T_144 = _T_142 | _T_143; // @[LZD.scala 49:16]
  assign _T_145 = ~ _T_143; // @[LZD.scala 49:27]
  assign _T_146 = _T_142 | _T_145; // @[LZD.scala 49:25]
  assign _T_147 = _T_80[2:0]; // @[LZD.scala 49:47]
  assign _T_148 = _T_141[2:0]; // @[LZD.scala 49:59]
  assign _T_149 = _T_142 ? _T_147 : _T_148; // @[LZD.scala 49:35]
  assign _T_151 = {_T_144,_T_146,_T_149}; // @[Cat.scala 29:58]
  assign _T_152 = _T_18[11:0]; // @[LZD.scala 44:32]
  assign _T_153 = _T_152[11:4]; // @[LZD.scala 43:32]
  assign _T_154 = _T_153[7:4]; // @[LZD.scala 43:32]
  assign _T_155 = _T_154[3:2]; // @[LZD.scala 43:32]
  assign _T_156 = _T_155 != 2'h0; // @[LZD.scala 39:14]
  assign _T_157 = _T_155[1]; // @[LZD.scala 39:21]
  assign _T_158 = _T_155[0]; // @[LZD.scala 39:30]
  assign _T_159 = ~ _T_158; // @[LZD.scala 39:27]
  assign _T_160 = _T_157 | _T_159; // @[LZD.scala 39:25]
  assign _T_161 = {_T_156,_T_160}; // @[Cat.scala 29:58]
  assign _T_162 = _T_154[1:0]; // @[LZD.scala 44:32]
  assign _T_163 = _T_162 != 2'h0; // @[LZD.scala 39:14]
  assign _T_164 = _T_162[1]; // @[LZD.scala 39:21]
  assign _T_165 = _T_162[0]; // @[LZD.scala 39:30]
  assign _T_166 = ~ _T_165; // @[LZD.scala 39:27]
  assign _T_167 = _T_164 | _T_166; // @[LZD.scala 39:25]
  assign _T_168 = {_T_163,_T_167}; // @[Cat.scala 29:58]
  assign _T_169 = _T_161[1]; // @[Shift.scala 12:21]
  assign _T_170 = _T_168[1]; // @[Shift.scala 12:21]
  assign _T_171 = _T_169 | _T_170; // @[LZD.scala 49:16]
  assign _T_172 = ~ _T_170; // @[LZD.scala 49:27]
  assign _T_173 = _T_169 | _T_172; // @[LZD.scala 49:25]
  assign _T_174 = _T_161[0:0]; // @[LZD.scala 49:47]
  assign _T_175 = _T_168[0:0]; // @[LZD.scala 49:59]
  assign _T_176 = _T_169 ? _T_174 : _T_175; // @[LZD.scala 49:35]
  assign _T_178 = {_T_171,_T_173,_T_176}; // @[Cat.scala 29:58]
  assign _T_179 = _T_153[3:0]; // @[LZD.scala 44:32]
  assign _T_180 = _T_179[3:2]; // @[LZD.scala 43:32]
  assign _T_181 = _T_180 != 2'h0; // @[LZD.scala 39:14]
  assign _T_182 = _T_180[1]; // @[LZD.scala 39:21]
  assign _T_183 = _T_180[0]; // @[LZD.scala 39:30]
  assign _T_184 = ~ _T_183; // @[LZD.scala 39:27]
  assign _T_185 = _T_182 | _T_184; // @[LZD.scala 39:25]
  assign _T_186 = {_T_181,_T_185}; // @[Cat.scala 29:58]
  assign _T_187 = _T_179[1:0]; // @[LZD.scala 44:32]
  assign _T_188 = _T_187 != 2'h0; // @[LZD.scala 39:14]
  assign _T_189 = _T_187[1]; // @[LZD.scala 39:21]
  assign _T_190 = _T_187[0]; // @[LZD.scala 39:30]
  assign _T_191 = ~ _T_190; // @[LZD.scala 39:27]
  assign _T_192 = _T_189 | _T_191; // @[LZD.scala 39:25]
  assign _T_193 = {_T_188,_T_192}; // @[Cat.scala 29:58]
  assign _T_194 = _T_186[1]; // @[Shift.scala 12:21]
  assign _T_195 = _T_193[1]; // @[Shift.scala 12:21]
  assign _T_196 = _T_194 | _T_195; // @[LZD.scala 49:16]
  assign _T_197 = ~ _T_195; // @[LZD.scala 49:27]
  assign _T_198 = _T_194 | _T_197; // @[LZD.scala 49:25]
  assign _T_199 = _T_186[0:0]; // @[LZD.scala 49:47]
  assign _T_200 = _T_193[0:0]; // @[LZD.scala 49:59]
  assign _T_201 = _T_194 ? _T_199 : _T_200; // @[LZD.scala 49:35]
  assign _T_203 = {_T_196,_T_198,_T_201}; // @[Cat.scala 29:58]
  assign _T_204 = _T_178[2]; // @[Shift.scala 12:21]
  assign _T_205 = _T_203[2]; // @[Shift.scala 12:21]
  assign _T_206 = _T_204 | _T_205; // @[LZD.scala 49:16]
  assign _T_207 = ~ _T_205; // @[LZD.scala 49:27]
  assign _T_208 = _T_204 | _T_207; // @[LZD.scala 49:25]
  assign _T_209 = _T_178[1:0]; // @[LZD.scala 49:47]
  assign _T_210 = _T_203[1:0]; // @[LZD.scala 49:59]
  assign _T_211 = _T_204 ? _T_209 : _T_210; // @[LZD.scala 49:35]
  assign _T_213 = {_T_206,_T_208,_T_211}; // @[Cat.scala 29:58]
  assign _T_214 = _T_152[3:0]; // @[LZD.scala 44:32]
  assign _T_215 = _T_214[3:2]; // @[LZD.scala 43:32]
  assign _T_216 = _T_215 != 2'h0; // @[LZD.scala 39:14]
  assign _T_217 = _T_215[1]; // @[LZD.scala 39:21]
  assign _T_218 = _T_215[0]; // @[LZD.scala 39:30]
  assign _T_219 = ~ _T_218; // @[LZD.scala 39:27]
  assign _T_220 = _T_217 | _T_219; // @[LZD.scala 39:25]
  assign _T_221 = {_T_216,_T_220}; // @[Cat.scala 29:58]
  assign _T_222 = _T_214[1:0]; // @[LZD.scala 44:32]
  assign _T_223 = _T_222 != 2'h0; // @[LZD.scala 39:14]
  assign _T_224 = _T_222[1]; // @[LZD.scala 39:21]
  assign _T_225 = _T_222[0]; // @[LZD.scala 39:30]
  assign _T_226 = ~ _T_225; // @[LZD.scala 39:27]
  assign _T_227 = _T_224 | _T_226; // @[LZD.scala 39:25]
  assign _T_228 = {_T_223,_T_227}; // @[Cat.scala 29:58]
  assign _T_229 = _T_221[1]; // @[Shift.scala 12:21]
  assign _T_230 = _T_228[1]; // @[Shift.scala 12:21]
  assign _T_231 = _T_229 | _T_230; // @[LZD.scala 49:16]
  assign _T_232 = ~ _T_230; // @[LZD.scala 49:27]
  assign _T_233 = _T_229 | _T_232; // @[LZD.scala 49:25]
  assign _T_234 = _T_221[0:0]; // @[LZD.scala 49:47]
  assign _T_235 = _T_228[0:0]; // @[LZD.scala 49:59]
  assign _T_236 = _T_229 ? _T_234 : _T_235; // @[LZD.scala 49:35]
  assign _T_238 = {_T_231,_T_233,_T_236}; // @[Cat.scala 29:58]
  assign _T_239 = _T_213[3]; // @[Shift.scala 12:21]
  assign _T_241 = _T_213[2:0]; // @[LZD.scala 55:32]
  assign _T_242 = _T_239 ? _T_241 : _T_238; // @[LZD.scala 55:20]
  assign _T_243 = {_T_239,_T_242}; // @[Cat.scala 29:58]
  assign _T_244 = _T_151[4]; // @[Shift.scala 12:21]
  assign _T_246 = _T_151[3:0]; // @[LZD.scala 55:32]
  assign _T_247 = _T_244 ? _T_246 : _T_243; // @[LZD.scala 55:20]
  assign _T_248 = {_T_244,_T_247}; // @[Cat.scala 29:58]
  assign _T_249 = ~ _T_248; // @[convert.scala 21:22]
  assign _T_250 = realA[26:0]; // @[convert.scala 22:36]
  assign _T_251 = _T_249 < 5'h1b; // @[Shift.scala 16:24]
  assign _T_253 = _T_249[4]; // @[Shift.scala 12:21]
  assign _T_254 = _T_250[10:0]; // @[Shift.scala 64:52]
  assign _T_256 = {_T_254,16'h0}; // @[Cat.scala 29:58]
  assign _T_257 = _T_253 ? _T_256 : _T_250; // @[Shift.scala 64:27]
  assign _T_258 = _T_249[3:0]; // @[Shift.scala 66:70]
  assign _T_259 = _T_258[3]; // @[Shift.scala 12:21]
  assign _T_260 = _T_257[18:0]; // @[Shift.scala 64:52]
  assign _T_262 = {_T_260,8'h0}; // @[Cat.scala 29:58]
  assign _T_263 = _T_259 ? _T_262 : _T_257; // @[Shift.scala 64:27]
  assign _T_264 = _T_258[2:0]; // @[Shift.scala 66:70]
  assign _T_265 = _T_264[2]; // @[Shift.scala 12:21]
  assign _T_266 = _T_263[22:0]; // @[Shift.scala 64:52]
  assign _T_268 = {_T_266,4'h0}; // @[Cat.scala 29:58]
  assign _T_269 = _T_265 ? _T_268 : _T_263; // @[Shift.scala 64:27]
  assign _T_270 = _T_264[1:0]; // @[Shift.scala 66:70]
  assign _T_271 = _T_270[1]; // @[Shift.scala 12:21]
  assign _T_272 = _T_269[24:0]; // @[Shift.scala 64:52]
  assign _T_274 = {_T_272,2'h0}; // @[Cat.scala 29:58]
  assign _T_275 = _T_271 ? _T_274 : _T_269; // @[Shift.scala 64:27]
  assign _T_276 = _T_270[0:0]; // @[Shift.scala 66:70]
  assign _T_278 = _T_275[25:0]; // @[Shift.scala 64:52]
  assign _T_279 = {_T_278,1'h0}; // @[Cat.scala 29:58]
  assign _T_280 = _T_276 ? _T_279 : _T_275; // @[Shift.scala 64:27]
  assign _T_281 = _T_251 ? _T_280 : 27'h0; // @[Shift.scala 16:10]
  assign _T_282 = _T_281[26:24]; // @[convert.scala 23:34]
  assign decA_fraction = _T_281[23:0]; // @[convert.scala 24:34]
  assign _T_284 = _T_15 == 1'h0; // @[convert.scala 25:26]
  assign _T_286 = _T_15 ? _T_249 : _T_248; // @[convert.scala 25:42]
  assign _T_289 = ~ _T_282; // @[convert.scala 26:67]
  assign _T_290 = _T_13 ? _T_289 : _T_282; // @[convert.scala 26:51]
  assign _T_291 = {_T_284,_T_286,_T_290}; // @[Cat.scala 29:58]
  assign _T_293 = realA[28:0]; // @[convert.scala 29:56]
  assign _T_294 = _T_293 != 29'h0; // @[convert.scala 29:60]
  assign _T_295 = ~ _T_294; // @[convert.scala 29:41]
  assign decA_isNaR = _T_13 & _T_295; // @[convert.scala 29:39]
  assign _T_298 = _T_13 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_298 & _T_295; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_291); // @[convert.scala 32:24]
  assign _T_307 = io_B[29]; // @[convert.scala 18:24]
  assign _T_308 = io_B[28]; // @[convert.scala 18:40]
  assign _T_309 = _T_307 ^ _T_308; // @[convert.scala 18:36]
  assign _T_310 = io_B[28:1]; // @[convert.scala 19:24]
  assign _T_311 = io_B[27:0]; // @[convert.scala 19:43]
  assign _T_312 = _T_310 ^ _T_311; // @[convert.scala 19:39]
  assign _T_313 = _T_312[27:12]; // @[LZD.scala 43:32]
  assign _T_314 = _T_313[15:8]; // @[LZD.scala 43:32]
  assign _T_315 = _T_314[7:4]; // @[LZD.scala 43:32]
  assign _T_316 = _T_315[3:2]; // @[LZD.scala 43:32]
  assign _T_317 = _T_316 != 2'h0; // @[LZD.scala 39:14]
  assign _T_318 = _T_316[1]; // @[LZD.scala 39:21]
  assign _T_319 = _T_316[0]; // @[LZD.scala 39:30]
  assign _T_320 = ~ _T_319; // @[LZD.scala 39:27]
  assign _T_321 = _T_318 | _T_320; // @[LZD.scala 39:25]
  assign _T_322 = {_T_317,_T_321}; // @[Cat.scala 29:58]
  assign _T_323 = _T_315[1:0]; // @[LZD.scala 44:32]
  assign _T_324 = _T_323 != 2'h0; // @[LZD.scala 39:14]
  assign _T_325 = _T_323[1]; // @[LZD.scala 39:21]
  assign _T_326 = _T_323[0]; // @[LZD.scala 39:30]
  assign _T_327 = ~ _T_326; // @[LZD.scala 39:27]
  assign _T_328 = _T_325 | _T_327; // @[LZD.scala 39:25]
  assign _T_329 = {_T_324,_T_328}; // @[Cat.scala 29:58]
  assign _T_330 = _T_322[1]; // @[Shift.scala 12:21]
  assign _T_331 = _T_329[1]; // @[Shift.scala 12:21]
  assign _T_332 = _T_330 | _T_331; // @[LZD.scala 49:16]
  assign _T_333 = ~ _T_331; // @[LZD.scala 49:27]
  assign _T_334 = _T_330 | _T_333; // @[LZD.scala 49:25]
  assign _T_335 = _T_322[0:0]; // @[LZD.scala 49:47]
  assign _T_336 = _T_329[0:0]; // @[LZD.scala 49:59]
  assign _T_337 = _T_330 ? _T_335 : _T_336; // @[LZD.scala 49:35]
  assign _T_339 = {_T_332,_T_334,_T_337}; // @[Cat.scala 29:58]
  assign _T_340 = _T_314[3:0]; // @[LZD.scala 44:32]
  assign _T_341 = _T_340[3:2]; // @[LZD.scala 43:32]
  assign _T_342 = _T_341 != 2'h0; // @[LZD.scala 39:14]
  assign _T_343 = _T_341[1]; // @[LZD.scala 39:21]
  assign _T_344 = _T_341[0]; // @[LZD.scala 39:30]
  assign _T_345 = ~ _T_344; // @[LZD.scala 39:27]
  assign _T_346 = _T_343 | _T_345; // @[LZD.scala 39:25]
  assign _T_347 = {_T_342,_T_346}; // @[Cat.scala 29:58]
  assign _T_348 = _T_340[1:0]; // @[LZD.scala 44:32]
  assign _T_349 = _T_348 != 2'h0; // @[LZD.scala 39:14]
  assign _T_350 = _T_348[1]; // @[LZD.scala 39:21]
  assign _T_351 = _T_348[0]; // @[LZD.scala 39:30]
  assign _T_352 = ~ _T_351; // @[LZD.scala 39:27]
  assign _T_353 = _T_350 | _T_352; // @[LZD.scala 39:25]
  assign _T_354 = {_T_349,_T_353}; // @[Cat.scala 29:58]
  assign _T_355 = _T_347[1]; // @[Shift.scala 12:21]
  assign _T_356 = _T_354[1]; // @[Shift.scala 12:21]
  assign _T_357 = _T_355 | _T_356; // @[LZD.scala 49:16]
  assign _T_358 = ~ _T_356; // @[LZD.scala 49:27]
  assign _T_359 = _T_355 | _T_358; // @[LZD.scala 49:25]
  assign _T_360 = _T_347[0:0]; // @[LZD.scala 49:47]
  assign _T_361 = _T_354[0:0]; // @[LZD.scala 49:59]
  assign _T_362 = _T_355 ? _T_360 : _T_361; // @[LZD.scala 49:35]
  assign _T_364 = {_T_357,_T_359,_T_362}; // @[Cat.scala 29:58]
  assign _T_365 = _T_339[2]; // @[Shift.scala 12:21]
  assign _T_366 = _T_364[2]; // @[Shift.scala 12:21]
  assign _T_367 = _T_365 | _T_366; // @[LZD.scala 49:16]
  assign _T_368 = ~ _T_366; // @[LZD.scala 49:27]
  assign _T_369 = _T_365 | _T_368; // @[LZD.scala 49:25]
  assign _T_370 = _T_339[1:0]; // @[LZD.scala 49:47]
  assign _T_371 = _T_364[1:0]; // @[LZD.scala 49:59]
  assign _T_372 = _T_365 ? _T_370 : _T_371; // @[LZD.scala 49:35]
  assign _T_374 = {_T_367,_T_369,_T_372}; // @[Cat.scala 29:58]
  assign _T_375 = _T_313[7:0]; // @[LZD.scala 44:32]
  assign _T_376 = _T_375[7:4]; // @[LZD.scala 43:32]
  assign _T_377 = _T_376[3:2]; // @[LZD.scala 43:32]
  assign _T_378 = _T_377 != 2'h0; // @[LZD.scala 39:14]
  assign _T_379 = _T_377[1]; // @[LZD.scala 39:21]
  assign _T_380 = _T_377[0]; // @[LZD.scala 39:30]
  assign _T_381 = ~ _T_380; // @[LZD.scala 39:27]
  assign _T_382 = _T_379 | _T_381; // @[LZD.scala 39:25]
  assign _T_383 = {_T_378,_T_382}; // @[Cat.scala 29:58]
  assign _T_384 = _T_376[1:0]; // @[LZD.scala 44:32]
  assign _T_385 = _T_384 != 2'h0; // @[LZD.scala 39:14]
  assign _T_386 = _T_384[1]; // @[LZD.scala 39:21]
  assign _T_387 = _T_384[0]; // @[LZD.scala 39:30]
  assign _T_388 = ~ _T_387; // @[LZD.scala 39:27]
  assign _T_389 = _T_386 | _T_388; // @[LZD.scala 39:25]
  assign _T_390 = {_T_385,_T_389}; // @[Cat.scala 29:58]
  assign _T_391 = _T_383[1]; // @[Shift.scala 12:21]
  assign _T_392 = _T_390[1]; // @[Shift.scala 12:21]
  assign _T_393 = _T_391 | _T_392; // @[LZD.scala 49:16]
  assign _T_394 = ~ _T_392; // @[LZD.scala 49:27]
  assign _T_395 = _T_391 | _T_394; // @[LZD.scala 49:25]
  assign _T_396 = _T_383[0:0]; // @[LZD.scala 49:47]
  assign _T_397 = _T_390[0:0]; // @[LZD.scala 49:59]
  assign _T_398 = _T_391 ? _T_396 : _T_397; // @[LZD.scala 49:35]
  assign _T_400 = {_T_393,_T_395,_T_398}; // @[Cat.scala 29:58]
  assign _T_401 = _T_375[3:0]; // @[LZD.scala 44:32]
  assign _T_402 = _T_401[3:2]; // @[LZD.scala 43:32]
  assign _T_403 = _T_402 != 2'h0; // @[LZD.scala 39:14]
  assign _T_404 = _T_402[1]; // @[LZD.scala 39:21]
  assign _T_405 = _T_402[0]; // @[LZD.scala 39:30]
  assign _T_406 = ~ _T_405; // @[LZD.scala 39:27]
  assign _T_407 = _T_404 | _T_406; // @[LZD.scala 39:25]
  assign _T_408 = {_T_403,_T_407}; // @[Cat.scala 29:58]
  assign _T_409 = _T_401[1:0]; // @[LZD.scala 44:32]
  assign _T_410 = _T_409 != 2'h0; // @[LZD.scala 39:14]
  assign _T_411 = _T_409[1]; // @[LZD.scala 39:21]
  assign _T_412 = _T_409[0]; // @[LZD.scala 39:30]
  assign _T_413 = ~ _T_412; // @[LZD.scala 39:27]
  assign _T_414 = _T_411 | _T_413; // @[LZD.scala 39:25]
  assign _T_415 = {_T_410,_T_414}; // @[Cat.scala 29:58]
  assign _T_416 = _T_408[1]; // @[Shift.scala 12:21]
  assign _T_417 = _T_415[1]; // @[Shift.scala 12:21]
  assign _T_418 = _T_416 | _T_417; // @[LZD.scala 49:16]
  assign _T_419 = ~ _T_417; // @[LZD.scala 49:27]
  assign _T_420 = _T_416 | _T_419; // @[LZD.scala 49:25]
  assign _T_421 = _T_408[0:0]; // @[LZD.scala 49:47]
  assign _T_422 = _T_415[0:0]; // @[LZD.scala 49:59]
  assign _T_423 = _T_416 ? _T_421 : _T_422; // @[LZD.scala 49:35]
  assign _T_425 = {_T_418,_T_420,_T_423}; // @[Cat.scala 29:58]
  assign _T_426 = _T_400[2]; // @[Shift.scala 12:21]
  assign _T_427 = _T_425[2]; // @[Shift.scala 12:21]
  assign _T_428 = _T_426 | _T_427; // @[LZD.scala 49:16]
  assign _T_429 = ~ _T_427; // @[LZD.scala 49:27]
  assign _T_430 = _T_426 | _T_429; // @[LZD.scala 49:25]
  assign _T_431 = _T_400[1:0]; // @[LZD.scala 49:47]
  assign _T_432 = _T_425[1:0]; // @[LZD.scala 49:59]
  assign _T_433 = _T_426 ? _T_431 : _T_432; // @[LZD.scala 49:35]
  assign _T_435 = {_T_428,_T_430,_T_433}; // @[Cat.scala 29:58]
  assign _T_436 = _T_374[3]; // @[Shift.scala 12:21]
  assign _T_437 = _T_435[3]; // @[Shift.scala 12:21]
  assign _T_438 = _T_436 | _T_437; // @[LZD.scala 49:16]
  assign _T_439 = ~ _T_437; // @[LZD.scala 49:27]
  assign _T_440 = _T_436 | _T_439; // @[LZD.scala 49:25]
  assign _T_441 = _T_374[2:0]; // @[LZD.scala 49:47]
  assign _T_442 = _T_435[2:0]; // @[LZD.scala 49:59]
  assign _T_443 = _T_436 ? _T_441 : _T_442; // @[LZD.scala 49:35]
  assign _T_445 = {_T_438,_T_440,_T_443}; // @[Cat.scala 29:58]
  assign _T_446 = _T_312[11:0]; // @[LZD.scala 44:32]
  assign _T_447 = _T_446[11:4]; // @[LZD.scala 43:32]
  assign _T_448 = _T_447[7:4]; // @[LZD.scala 43:32]
  assign _T_449 = _T_448[3:2]; // @[LZD.scala 43:32]
  assign _T_450 = _T_449 != 2'h0; // @[LZD.scala 39:14]
  assign _T_451 = _T_449[1]; // @[LZD.scala 39:21]
  assign _T_452 = _T_449[0]; // @[LZD.scala 39:30]
  assign _T_453 = ~ _T_452; // @[LZD.scala 39:27]
  assign _T_454 = _T_451 | _T_453; // @[LZD.scala 39:25]
  assign _T_455 = {_T_450,_T_454}; // @[Cat.scala 29:58]
  assign _T_456 = _T_448[1:0]; // @[LZD.scala 44:32]
  assign _T_457 = _T_456 != 2'h0; // @[LZD.scala 39:14]
  assign _T_458 = _T_456[1]; // @[LZD.scala 39:21]
  assign _T_459 = _T_456[0]; // @[LZD.scala 39:30]
  assign _T_460 = ~ _T_459; // @[LZD.scala 39:27]
  assign _T_461 = _T_458 | _T_460; // @[LZD.scala 39:25]
  assign _T_462 = {_T_457,_T_461}; // @[Cat.scala 29:58]
  assign _T_463 = _T_455[1]; // @[Shift.scala 12:21]
  assign _T_464 = _T_462[1]; // @[Shift.scala 12:21]
  assign _T_465 = _T_463 | _T_464; // @[LZD.scala 49:16]
  assign _T_466 = ~ _T_464; // @[LZD.scala 49:27]
  assign _T_467 = _T_463 | _T_466; // @[LZD.scala 49:25]
  assign _T_468 = _T_455[0:0]; // @[LZD.scala 49:47]
  assign _T_469 = _T_462[0:0]; // @[LZD.scala 49:59]
  assign _T_470 = _T_463 ? _T_468 : _T_469; // @[LZD.scala 49:35]
  assign _T_472 = {_T_465,_T_467,_T_470}; // @[Cat.scala 29:58]
  assign _T_473 = _T_447[3:0]; // @[LZD.scala 44:32]
  assign _T_474 = _T_473[3:2]; // @[LZD.scala 43:32]
  assign _T_475 = _T_474 != 2'h0; // @[LZD.scala 39:14]
  assign _T_476 = _T_474[1]; // @[LZD.scala 39:21]
  assign _T_477 = _T_474[0]; // @[LZD.scala 39:30]
  assign _T_478 = ~ _T_477; // @[LZD.scala 39:27]
  assign _T_479 = _T_476 | _T_478; // @[LZD.scala 39:25]
  assign _T_480 = {_T_475,_T_479}; // @[Cat.scala 29:58]
  assign _T_481 = _T_473[1:0]; // @[LZD.scala 44:32]
  assign _T_482 = _T_481 != 2'h0; // @[LZD.scala 39:14]
  assign _T_483 = _T_481[1]; // @[LZD.scala 39:21]
  assign _T_484 = _T_481[0]; // @[LZD.scala 39:30]
  assign _T_485 = ~ _T_484; // @[LZD.scala 39:27]
  assign _T_486 = _T_483 | _T_485; // @[LZD.scala 39:25]
  assign _T_487 = {_T_482,_T_486}; // @[Cat.scala 29:58]
  assign _T_488 = _T_480[1]; // @[Shift.scala 12:21]
  assign _T_489 = _T_487[1]; // @[Shift.scala 12:21]
  assign _T_490 = _T_488 | _T_489; // @[LZD.scala 49:16]
  assign _T_491 = ~ _T_489; // @[LZD.scala 49:27]
  assign _T_492 = _T_488 | _T_491; // @[LZD.scala 49:25]
  assign _T_493 = _T_480[0:0]; // @[LZD.scala 49:47]
  assign _T_494 = _T_487[0:0]; // @[LZD.scala 49:59]
  assign _T_495 = _T_488 ? _T_493 : _T_494; // @[LZD.scala 49:35]
  assign _T_497 = {_T_490,_T_492,_T_495}; // @[Cat.scala 29:58]
  assign _T_498 = _T_472[2]; // @[Shift.scala 12:21]
  assign _T_499 = _T_497[2]; // @[Shift.scala 12:21]
  assign _T_500 = _T_498 | _T_499; // @[LZD.scala 49:16]
  assign _T_501 = ~ _T_499; // @[LZD.scala 49:27]
  assign _T_502 = _T_498 | _T_501; // @[LZD.scala 49:25]
  assign _T_503 = _T_472[1:0]; // @[LZD.scala 49:47]
  assign _T_504 = _T_497[1:0]; // @[LZD.scala 49:59]
  assign _T_505 = _T_498 ? _T_503 : _T_504; // @[LZD.scala 49:35]
  assign _T_507 = {_T_500,_T_502,_T_505}; // @[Cat.scala 29:58]
  assign _T_508 = _T_446[3:0]; // @[LZD.scala 44:32]
  assign _T_509 = _T_508[3:2]; // @[LZD.scala 43:32]
  assign _T_510 = _T_509 != 2'h0; // @[LZD.scala 39:14]
  assign _T_511 = _T_509[1]; // @[LZD.scala 39:21]
  assign _T_512 = _T_509[0]; // @[LZD.scala 39:30]
  assign _T_513 = ~ _T_512; // @[LZD.scala 39:27]
  assign _T_514 = _T_511 | _T_513; // @[LZD.scala 39:25]
  assign _T_515 = {_T_510,_T_514}; // @[Cat.scala 29:58]
  assign _T_516 = _T_508[1:0]; // @[LZD.scala 44:32]
  assign _T_517 = _T_516 != 2'h0; // @[LZD.scala 39:14]
  assign _T_518 = _T_516[1]; // @[LZD.scala 39:21]
  assign _T_519 = _T_516[0]; // @[LZD.scala 39:30]
  assign _T_520 = ~ _T_519; // @[LZD.scala 39:27]
  assign _T_521 = _T_518 | _T_520; // @[LZD.scala 39:25]
  assign _T_522 = {_T_517,_T_521}; // @[Cat.scala 29:58]
  assign _T_523 = _T_515[1]; // @[Shift.scala 12:21]
  assign _T_524 = _T_522[1]; // @[Shift.scala 12:21]
  assign _T_525 = _T_523 | _T_524; // @[LZD.scala 49:16]
  assign _T_526 = ~ _T_524; // @[LZD.scala 49:27]
  assign _T_527 = _T_523 | _T_526; // @[LZD.scala 49:25]
  assign _T_528 = _T_515[0:0]; // @[LZD.scala 49:47]
  assign _T_529 = _T_522[0:0]; // @[LZD.scala 49:59]
  assign _T_530 = _T_523 ? _T_528 : _T_529; // @[LZD.scala 49:35]
  assign _T_532 = {_T_525,_T_527,_T_530}; // @[Cat.scala 29:58]
  assign _T_533 = _T_507[3]; // @[Shift.scala 12:21]
  assign _T_535 = _T_507[2:0]; // @[LZD.scala 55:32]
  assign _T_536 = _T_533 ? _T_535 : _T_532; // @[LZD.scala 55:20]
  assign _T_537 = {_T_533,_T_536}; // @[Cat.scala 29:58]
  assign _T_538 = _T_445[4]; // @[Shift.scala 12:21]
  assign _T_540 = _T_445[3:0]; // @[LZD.scala 55:32]
  assign _T_541 = _T_538 ? _T_540 : _T_537; // @[LZD.scala 55:20]
  assign _T_542 = {_T_538,_T_541}; // @[Cat.scala 29:58]
  assign _T_543 = ~ _T_542; // @[convert.scala 21:22]
  assign _T_544 = io_B[26:0]; // @[convert.scala 22:36]
  assign _T_545 = _T_543 < 5'h1b; // @[Shift.scala 16:24]
  assign _T_547 = _T_543[4]; // @[Shift.scala 12:21]
  assign _T_548 = _T_544[10:0]; // @[Shift.scala 64:52]
  assign _T_550 = {_T_548,16'h0}; // @[Cat.scala 29:58]
  assign _T_551 = _T_547 ? _T_550 : _T_544; // @[Shift.scala 64:27]
  assign _T_552 = _T_543[3:0]; // @[Shift.scala 66:70]
  assign _T_553 = _T_552[3]; // @[Shift.scala 12:21]
  assign _T_554 = _T_551[18:0]; // @[Shift.scala 64:52]
  assign _T_556 = {_T_554,8'h0}; // @[Cat.scala 29:58]
  assign _T_557 = _T_553 ? _T_556 : _T_551; // @[Shift.scala 64:27]
  assign _T_558 = _T_552[2:0]; // @[Shift.scala 66:70]
  assign _T_559 = _T_558[2]; // @[Shift.scala 12:21]
  assign _T_560 = _T_557[22:0]; // @[Shift.scala 64:52]
  assign _T_562 = {_T_560,4'h0}; // @[Cat.scala 29:58]
  assign _T_563 = _T_559 ? _T_562 : _T_557; // @[Shift.scala 64:27]
  assign _T_564 = _T_558[1:0]; // @[Shift.scala 66:70]
  assign _T_565 = _T_564[1]; // @[Shift.scala 12:21]
  assign _T_566 = _T_563[24:0]; // @[Shift.scala 64:52]
  assign _T_568 = {_T_566,2'h0}; // @[Cat.scala 29:58]
  assign _T_569 = _T_565 ? _T_568 : _T_563; // @[Shift.scala 64:27]
  assign _T_570 = _T_564[0:0]; // @[Shift.scala 66:70]
  assign _T_572 = _T_569[25:0]; // @[Shift.scala 64:52]
  assign _T_573 = {_T_572,1'h0}; // @[Cat.scala 29:58]
  assign _T_574 = _T_570 ? _T_573 : _T_569; // @[Shift.scala 64:27]
  assign _T_575 = _T_545 ? _T_574 : 27'h0; // @[Shift.scala 16:10]
  assign _T_576 = _T_575[26:24]; // @[convert.scala 23:34]
  assign decB_fraction = _T_575[23:0]; // @[convert.scala 24:34]
  assign _T_578 = _T_309 == 1'h0; // @[convert.scala 25:26]
  assign _T_580 = _T_309 ? _T_543 : _T_542; // @[convert.scala 25:42]
  assign _T_583 = ~ _T_576; // @[convert.scala 26:67]
  assign _T_584 = _T_307 ? _T_583 : _T_576; // @[convert.scala 26:51]
  assign _T_585 = {_T_578,_T_580,_T_584}; // @[Cat.scala 29:58]
  assign _T_587 = io_B[28:0]; // @[convert.scala 29:56]
  assign _T_588 = _T_587 != 29'h0; // @[convert.scala 29:60]
  assign _T_589 = ~ _T_588; // @[convert.scala 29:41]
  assign decB_isNaR = _T_307 & _T_589; // @[convert.scala 29:39]
  assign _T_592 = _T_307 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_592 & _T_589; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_585); // @[convert.scala 32:24]
  assign _T_601 = realC[29]; // @[convert.scala 18:24]
  assign _T_602 = realC[28]; // @[convert.scala 18:40]
  assign _T_603 = _T_601 ^ _T_602; // @[convert.scala 18:36]
  assign _T_604 = realC[28:1]; // @[convert.scala 19:24]
  assign _T_605 = realC[27:0]; // @[convert.scala 19:43]
  assign _T_606 = _T_604 ^ _T_605; // @[convert.scala 19:39]
  assign _T_607 = _T_606[27:12]; // @[LZD.scala 43:32]
  assign _T_608 = _T_607[15:8]; // @[LZD.scala 43:32]
  assign _T_609 = _T_608[7:4]; // @[LZD.scala 43:32]
  assign _T_610 = _T_609[3:2]; // @[LZD.scala 43:32]
  assign _T_611 = _T_610 != 2'h0; // @[LZD.scala 39:14]
  assign _T_612 = _T_610[1]; // @[LZD.scala 39:21]
  assign _T_613 = _T_610[0]; // @[LZD.scala 39:30]
  assign _T_614 = ~ _T_613; // @[LZD.scala 39:27]
  assign _T_615 = _T_612 | _T_614; // @[LZD.scala 39:25]
  assign _T_616 = {_T_611,_T_615}; // @[Cat.scala 29:58]
  assign _T_617 = _T_609[1:0]; // @[LZD.scala 44:32]
  assign _T_618 = _T_617 != 2'h0; // @[LZD.scala 39:14]
  assign _T_619 = _T_617[1]; // @[LZD.scala 39:21]
  assign _T_620 = _T_617[0]; // @[LZD.scala 39:30]
  assign _T_621 = ~ _T_620; // @[LZD.scala 39:27]
  assign _T_622 = _T_619 | _T_621; // @[LZD.scala 39:25]
  assign _T_623 = {_T_618,_T_622}; // @[Cat.scala 29:58]
  assign _T_624 = _T_616[1]; // @[Shift.scala 12:21]
  assign _T_625 = _T_623[1]; // @[Shift.scala 12:21]
  assign _T_626 = _T_624 | _T_625; // @[LZD.scala 49:16]
  assign _T_627 = ~ _T_625; // @[LZD.scala 49:27]
  assign _T_628 = _T_624 | _T_627; // @[LZD.scala 49:25]
  assign _T_629 = _T_616[0:0]; // @[LZD.scala 49:47]
  assign _T_630 = _T_623[0:0]; // @[LZD.scala 49:59]
  assign _T_631 = _T_624 ? _T_629 : _T_630; // @[LZD.scala 49:35]
  assign _T_633 = {_T_626,_T_628,_T_631}; // @[Cat.scala 29:58]
  assign _T_634 = _T_608[3:0]; // @[LZD.scala 44:32]
  assign _T_635 = _T_634[3:2]; // @[LZD.scala 43:32]
  assign _T_636 = _T_635 != 2'h0; // @[LZD.scala 39:14]
  assign _T_637 = _T_635[1]; // @[LZD.scala 39:21]
  assign _T_638 = _T_635[0]; // @[LZD.scala 39:30]
  assign _T_639 = ~ _T_638; // @[LZD.scala 39:27]
  assign _T_640 = _T_637 | _T_639; // @[LZD.scala 39:25]
  assign _T_641 = {_T_636,_T_640}; // @[Cat.scala 29:58]
  assign _T_642 = _T_634[1:0]; // @[LZD.scala 44:32]
  assign _T_643 = _T_642 != 2'h0; // @[LZD.scala 39:14]
  assign _T_644 = _T_642[1]; // @[LZD.scala 39:21]
  assign _T_645 = _T_642[0]; // @[LZD.scala 39:30]
  assign _T_646 = ~ _T_645; // @[LZD.scala 39:27]
  assign _T_647 = _T_644 | _T_646; // @[LZD.scala 39:25]
  assign _T_648 = {_T_643,_T_647}; // @[Cat.scala 29:58]
  assign _T_649 = _T_641[1]; // @[Shift.scala 12:21]
  assign _T_650 = _T_648[1]; // @[Shift.scala 12:21]
  assign _T_651 = _T_649 | _T_650; // @[LZD.scala 49:16]
  assign _T_652 = ~ _T_650; // @[LZD.scala 49:27]
  assign _T_653 = _T_649 | _T_652; // @[LZD.scala 49:25]
  assign _T_654 = _T_641[0:0]; // @[LZD.scala 49:47]
  assign _T_655 = _T_648[0:0]; // @[LZD.scala 49:59]
  assign _T_656 = _T_649 ? _T_654 : _T_655; // @[LZD.scala 49:35]
  assign _T_658 = {_T_651,_T_653,_T_656}; // @[Cat.scala 29:58]
  assign _T_659 = _T_633[2]; // @[Shift.scala 12:21]
  assign _T_660 = _T_658[2]; // @[Shift.scala 12:21]
  assign _T_661 = _T_659 | _T_660; // @[LZD.scala 49:16]
  assign _T_662 = ~ _T_660; // @[LZD.scala 49:27]
  assign _T_663 = _T_659 | _T_662; // @[LZD.scala 49:25]
  assign _T_664 = _T_633[1:0]; // @[LZD.scala 49:47]
  assign _T_665 = _T_658[1:0]; // @[LZD.scala 49:59]
  assign _T_666 = _T_659 ? _T_664 : _T_665; // @[LZD.scala 49:35]
  assign _T_668 = {_T_661,_T_663,_T_666}; // @[Cat.scala 29:58]
  assign _T_669 = _T_607[7:0]; // @[LZD.scala 44:32]
  assign _T_670 = _T_669[7:4]; // @[LZD.scala 43:32]
  assign _T_671 = _T_670[3:2]; // @[LZD.scala 43:32]
  assign _T_672 = _T_671 != 2'h0; // @[LZD.scala 39:14]
  assign _T_673 = _T_671[1]; // @[LZD.scala 39:21]
  assign _T_674 = _T_671[0]; // @[LZD.scala 39:30]
  assign _T_675 = ~ _T_674; // @[LZD.scala 39:27]
  assign _T_676 = _T_673 | _T_675; // @[LZD.scala 39:25]
  assign _T_677 = {_T_672,_T_676}; // @[Cat.scala 29:58]
  assign _T_678 = _T_670[1:0]; // @[LZD.scala 44:32]
  assign _T_679 = _T_678 != 2'h0; // @[LZD.scala 39:14]
  assign _T_680 = _T_678[1]; // @[LZD.scala 39:21]
  assign _T_681 = _T_678[0]; // @[LZD.scala 39:30]
  assign _T_682 = ~ _T_681; // @[LZD.scala 39:27]
  assign _T_683 = _T_680 | _T_682; // @[LZD.scala 39:25]
  assign _T_684 = {_T_679,_T_683}; // @[Cat.scala 29:58]
  assign _T_685 = _T_677[1]; // @[Shift.scala 12:21]
  assign _T_686 = _T_684[1]; // @[Shift.scala 12:21]
  assign _T_687 = _T_685 | _T_686; // @[LZD.scala 49:16]
  assign _T_688 = ~ _T_686; // @[LZD.scala 49:27]
  assign _T_689 = _T_685 | _T_688; // @[LZD.scala 49:25]
  assign _T_690 = _T_677[0:0]; // @[LZD.scala 49:47]
  assign _T_691 = _T_684[0:0]; // @[LZD.scala 49:59]
  assign _T_692 = _T_685 ? _T_690 : _T_691; // @[LZD.scala 49:35]
  assign _T_694 = {_T_687,_T_689,_T_692}; // @[Cat.scala 29:58]
  assign _T_695 = _T_669[3:0]; // @[LZD.scala 44:32]
  assign _T_696 = _T_695[3:2]; // @[LZD.scala 43:32]
  assign _T_697 = _T_696 != 2'h0; // @[LZD.scala 39:14]
  assign _T_698 = _T_696[1]; // @[LZD.scala 39:21]
  assign _T_699 = _T_696[0]; // @[LZD.scala 39:30]
  assign _T_700 = ~ _T_699; // @[LZD.scala 39:27]
  assign _T_701 = _T_698 | _T_700; // @[LZD.scala 39:25]
  assign _T_702 = {_T_697,_T_701}; // @[Cat.scala 29:58]
  assign _T_703 = _T_695[1:0]; // @[LZD.scala 44:32]
  assign _T_704 = _T_703 != 2'h0; // @[LZD.scala 39:14]
  assign _T_705 = _T_703[1]; // @[LZD.scala 39:21]
  assign _T_706 = _T_703[0]; // @[LZD.scala 39:30]
  assign _T_707 = ~ _T_706; // @[LZD.scala 39:27]
  assign _T_708 = _T_705 | _T_707; // @[LZD.scala 39:25]
  assign _T_709 = {_T_704,_T_708}; // @[Cat.scala 29:58]
  assign _T_710 = _T_702[1]; // @[Shift.scala 12:21]
  assign _T_711 = _T_709[1]; // @[Shift.scala 12:21]
  assign _T_712 = _T_710 | _T_711; // @[LZD.scala 49:16]
  assign _T_713 = ~ _T_711; // @[LZD.scala 49:27]
  assign _T_714 = _T_710 | _T_713; // @[LZD.scala 49:25]
  assign _T_715 = _T_702[0:0]; // @[LZD.scala 49:47]
  assign _T_716 = _T_709[0:0]; // @[LZD.scala 49:59]
  assign _T_717 = _T_710 ? _T_715 : _T_716; // @[LZD.scala 49:35]
  assign _T_719 = {_T_712,_T_714,_T_717}; // @[Cat.scala 29:58]
  assign _T_720 = _T_694[2]; // @[Shift.scala 12:21]
  assign _T_721 = _T_719[2]; // @[Shift.scala 12:21]
  assign _T_722 = _T_720 | _T_721; // @[LZD.scala 49:16]
  assign _T_723 = ~ _T_721; // @[LZD.scala 49:27]
  assign _T_724 = _T_720 | _T_723; // @[LZD.scala 49:25]
  assign _T_725 = _T_694[1:0]; // @[LZD.scala 49:47]
  assign _T_726 = _T_719[1:0]; // @[LZD.scala 49:59]
  assign _T_727 = _T_720 ? _T_725 : _T_726; // @[LZD.scala 49:35]
  assign _T_729 = {_T_722,_T_724,_T_727}; // @[Cat.scala 29:58]
  assign _T_730 = _T_668[3]; // @[Shift.scala 12:21]
  assign _T_731 = _T_729[3]; // @[Shift.scala 12:21]
  assign _T_732 = _T_730 | _T_731; // @[LZD.scala 49:16]
  assign _T_733 = ~ _T_731; // @[LZD.scala 49:27]
  assign _T_734 = _T_730 | _T_733; // @[LZD.scala 49:25]
  assign _T_735 = _T_668[2:0]; // @[LZD.scala 49:47]
  assign _T_736 = _T_729[2:0]; // @[LZD.scala 49:59]
  assign _T_737 = _T_730 ? _T_735 : _T_736; // @[LZD.scala 49:35]
  assign _T_739 = {_T_732,_T_734,_T_737}; // @[Cat.scala 29:58]
  assign _T_740 = _T_606[11:0]; // @[LZD.scala 44:32]
  assign _T_741 = _T_740[11:4]; // @[LZD.scala 43:32]
  assign _T_742 = _T_741[7:4]; // @[LZD.scala 43:32]
  assign _T_743 = _T_742[3:2]; // @[LZD.scala 43:32]
  assign _T_744 = _T_743 != 2'h0; // @[LZD.scala 39:14]
  assign _T_745 = _T_743[1]; // @[LZD.scala 39:21]
  assign _T_746 = _T_743[0]; // @[LZD.scala 39:30]
  assign _T_747 = ~ _T_746; // @[LZD.scala 39:27]
  assign _T_748 = _T_745 | _T_747; // @[LZD.scala 39:25]
  assign _T_749 = {_T_744,_T_748}; // @[Cat.scala 29:58]
  assign _T_750 = _T_742[1:0]; // @[LZD.scala 44:32]
  assign _T_751 = _T_750 != 2'h0; // @[LZD.scala 39:14]
  assign _T_752 = _T_750[1]; // @[LZD.scala 39:21]
  assign _T_753 = _T_750[0]; // @[LZD.scala 39:30]
  assign _T_754 = ~ _T_753; // @[LZD.scala 39:27]
  assign _T_755 = _T_752 | _T_754; // @[LZD.scala 39:25]
  assign _T_756 = {_T_751,_T_755}; // @[Cat.scala 29:58]
  assign _T_757 = _T_749[1]; // @[Shift.scala 12:21]
  assign _T_758 = _T_756[1]; // @[Shift.scala 12:21]
  assign _T_759 = _T_757 | _T_758; // @[LZD.scala 49:16]
  assign _T_760 = ~ _T_758; // @[LZD.scala 49:27]
  assign _T_761 = _T_757 | _T_760; // @[LZD.scala 49:25]
  assign _T_762 = _T_749[0:0]; // @[LZD.scala 49:47]
  assign _T_763 = _T_756[0:0]; // @[LZD.scala 49:59]
  assign _T_764 = _T_757 ? _T_762 : _T_763; // @[LZD.scala 49:35]
  assign _T_766 = {_T_759,_T_761,_T_764}; // @[Cat.scala 29:58]
  assign _T_767 = _T_741[3:0]; // @[LZD.scala 44:32]
  assign _T_768 = _T_767[3:2]; // @[LZD.scala 43:32]
  assign _T_769 = _T_768 != 2'h0; // @[LZD.scala 39:14]
  assign _T_770 = _T_768[1]; // @[LZD.scala 39:21]
  assign _T_771 = _T_768[0]; // @[LZD.scala 39:30]
  assign _T_772 = ~ _T_771; // @[LZD.scala 39:27]
  assign _T_773 = _T_770 | _T_772; // @[LZD.scala 39:25]
  assign _T_774 = {_T_769,_T_773}; // @[Cat.scala 29:58]
  assign _T_775 = _T_767[1:0]; // @[LZD.scala 44:32]
  assign _T_776 = _T_775 != 2'h0; // @[LZD.scala 39:14]
  assign _T_777 = _T_775[1]; // @[LZD.scala 39:21]
  assign _T_778 = _T_775[0]; // @[LZD.scala 39:30]
  assign _T_779 = ~ _T_778; // @[LZD.scala 39:27]
  assign _T_780 = _T_777 | _T_779; // @[LZD.scala 39:25]
  assign _T_781 = {_T_776,_T_780}; // @[Cat.scala 29:58]
  assign _T_782 = _T_774[1]; // @[Shift.scala 12:21]
  assign _T_783 = _T_781[1]; // @[Shift.scala 12:21]
  assign _T_784 = _T_782 | _T_783; // @[LZD.scala 49:16]
  assign _T_785 = ~ _T_783; // @[LZD.scala 49:27]
  assign _T_786 = _T_782 | _T_785; // @[LZD.scala 49:25]
  assign _T_787 = _T_774[0:0]; // @[LZD.scala 49:47]
  assign _T_788 = _T_781[0:0]; // @[LZD.scala 49:59]
  assign _T_789 = _T_782 ? _T_787 : _T_788; // @[LZD.scala 49:35]
  assign _T_791 = {_T_784,_T_786,_T_789}; // @[Cat.scala 29:58]
  assign _T_792 = _T_766[2]; // @[Shift.scala 12:21]
  assign _T_793 = _T_791[2]; // @[Shift.scala 12:21]
  assign _T_794 = _T_792 | _T_793; // @[LZD.scala 49:16]
  assign _T_795 = ~ _T_793; // @[LZD.scala 49:27]
  assign _T_796 = _T_792 | _T_795; // @[LZD.scala 49:25]
  assign _T_797 = _T_766[1:0]; // @[LZD.scala 49:47]
  assign _T_798 = _T_791[1:0]; // @[LZD.scala 49:59]
  assign _T_799 = _T_792 ? _T_797 : _T_798; // @[LZD.scala 49:35]
  assign _T_801 = {_T_794,_T_796,_T_799}; // @[Cat.scala 29:58]
  assign _T_802 = _T_740[3:0]; // @[LZD.scala 44:32]
  assign _T_803 = _T_802[3:2]; // @[LZD.scala 43:32]
  assign _T_804 = _T_803 != 2'h0; // @[LZD.scala 39:14]
  assign _T_805 = _T_803[1]; // @[LZD.scala 39:21]
  assign _T_806 = _T_803[0]; // @[LZD.scala 39:30]
  assign _T_807 = ~ _T_806; // @[LZD.scala 39:27]
  assign _T_808 = _T_805 | _T_807; // @[LZD.scala 39:25]
  assign _T_809 = {_T_804,_T_808}; // @[Cat.scala 29:58]
  assign _T_810 = _T_802[1:0]; // @[LZD.scala 44:32]
  assign _T_811 = _T_810 != 2'h0; // @[LZD.scala 39:14]
  assign _T_812 = _T_810[1]; // @[LZD.scala 39:21]
  assign _T_813 = _T_810[0]; // @[LZD.scala 39:30]
  assign _T_814 = ~ _T_813; // @[LZD.scala 39:27]
  assign _T_815 = _T_812 | _T_814; // @[LZD.scala 39:25]
  assign _T_816 = {_T_811,_T_815}; // @[Cat.scala 29:58]
  assign _T_817 = _T_809[1]; // @[Shift.scala 12:21]
  assign _T_818 = _T_816[1]; // @[Shift.scala 12:21]
  assign _T_819 = _T_817 | _T_818; // @[LZD.scala 49:16]
  assign _T_820 = ~ _T_818; // @[LZD.scala 49:27]
  assign _T_821 = _T_817 | _T_820; // @[LZD.scala 49:25]
  assign _T_822 = _T_809[0:0]; // @[LZD.scala 49:47]
  assign _T_823 = _T_816[0:0]; // @[LZD.scala 49:59]
  assign _T_824 = _T_817 ? _T_822 : _T_823; // @[LZD.scala 49:35]
  assign _T_826 = {_T_819,_T_821,_T_824}; // @[Cat.scala 29:58]
  assign _T_827 = _T_801[3]; // @[Shift.scala 12:21]
  assign _T_829 = _T_801[2:0]; // @[LZD.scala 55:32]
  assign _T_830 = _T_827 ? _T_829 : _T_826; // @[LZD.scala 55:20]
  assign _T_831 = {_T_827,_T_830}; // @[Cat.scala 29:58]
  assign _T_832 = _T_739[4]; // @[Shift.scala 12:21]
  assign _T_834 = _T_739[3:0]; // @[LZD.scala 55:32]
  assign _T_835 = _T_832 ? _T_834 : _T_831; // @[LZD.scala 55:20]
  assign _T_836 = {_T_832,_T_835}; // @[Cat.scala 29:58]
  assign _T_837 = ~ _T_836; // @[convert.scala 21:22]
  assign _T_838 = realC[26:0]; // @[convert.scala 22:36]
  assign _T_839 = _T_837 < 5'h1b; // @[Shift.scala 16:24]
  assign _T_841 = _T_837[4]; // @[Shift.scala 12:21]
  assign _T_842 = _T_838[10:0]; // @[Shift.scala 64:52]
  assign _T_844 = {_T_842,16'h0}; // @[Cat.scala 29:58]
  assign _T_845 = _T_841 ? _T_844 : _T_838; // @[Shift.scala 64:27]
  assign _T_846 = _T_837[3:0]; // @[Shift.scala 66:70]
  assign _T_847 = _T_846[3]; // @[Shift.scala 12:21]
  assign _T_848 = _T_845[18:0]; // @[Shift.scala 64:52]
  assign _T_850 = {_T_848,8'h0}; // @[Cat.scala 29:58]
  assign _T_851 = _T_847 ? _T_850 : _T_845; // @[Shift.scala 64:27]
  assign _T_852 = _T_846[2:0]; // @[Shift.scala 66:70]
  assign _T_853 = _T_852[2]; // @[Shift.scala 12:21]
  assign _T_854 = _T_851[22:0]; // @[Shift.scala 64:52]
  assign _T_856 = {_T_854,4'h0}; // @[Cat.scala 29:58]
  assign _T_857 = _T_853 ? _T_856 : _T_851; // @[Shift.scala 64:27]
  assign _T_858 = _T_852[1:0]; // @[Shift.scala 66:70]
  assign _T_859 = _T_858[1]; // @[Shift.scala 12:21]
  assign _T_860 = _T_857[24:0]; // @[Shift.scala 64:52]
  assign _T_862 = {_T_860,2'h0}; // @[Cat.scala 29:58]
  assign _T_863 = _T_859 ? _T_862 : _T_857; // @[Shift.scala 64:27]
  assign _T_864 = _T_858[0:0]; // @[Shift.scala 66:70]
  assign _T_866 = _T_863[25:0]; // @[Shift.scala 64:52]
  assign _T_867 = {_T_866,1'h0}; // @[Cat.scala 29:58]
  assign _T_868 = _T_864 ? _T_867 : _T_863; // @[Shift.scala 64:27]
  assign _T_869 = _T_839 ? _T_868 : 27'h0; // @[Shift.scala 16:10]
  assign _T_870 = _T_869[26:24]; // @[convert.scala 23:34]
  assign decC_fraction = _T_869[23:0]; // @[convert.scala 24:34]
  assign _T_872 = _T_603 == 1'h0; // @[convert.scala 25:26]
  assign _T_874 = _T_603 ? _T_837 : _T_836; // @[convert.scala 25:42]
  assign _T_877 = ~ _T_870; // @[convert.scala 26:67]
  assign _T_878 = _T_601 ? _T_877 : _T_870; // @[convert.scala 26:51]
  assign _T_879 = {_T_872,_T_874,_T_878}; // @[Cat.scala 29:58]
  assign _T_881 = realC[28:0]; // @[convert.scala 29:56]
  assign _T_882 = _T_881 != 29'h0; // @[convert.scala 29:60]
  assign _T_883 = ~ _T_882; // @[convert.scala 29:41]
  assign decC_isNaR = _T_601 & _T_883; // @[convert.scala 29:39]
  assign _T_886 = _T_601 == 1'h0; // @[convert.scala 30:19]
  assign decC_isZero = _T_886 & _T_883; // @[convert.scala 30:41]
  assign decC_scale = $signed(_T_879); // @[convert.scala 32:24]
  assign _T_894 = decA_isNaR | decB_isNaR; // @[PositFMA.scala 58:30]
  assign outIsNaR = _T_894 | decC_isNaR; // @[PositFMA.scala 58:44]
  assign _T_895 = ~ _T_13; // @[PositFMA.scala 59:34]
  assign _T_896 = ~ decA_isZero; // @[PositFMA.scala 59:47]
  assign _T_897 = _T_895 & _T_896; // @[PositFMA.scala 59:45]
  assign _T_899 = {_T_13,_T_897,decA_fraction}; // @[Cat.scala 29:58]
  assign sigA = $signed(_T_899); // @[PositFMA.scala 59:76]
  assign _T_900 = ~ _T_307; // @[PositFMA.scala 60:34]
  assign _T_901 = ~ decB_isZero; // @[PositFMA.scala 60:47]
  assign _T_902 = _T_900 & _T_901; // @[PositFMA.scala 60:45]
  assign _T_904 = {_T_307,_T_902,decB_fraction}; // @[Cat.scala 29:58]
  assign sigB = $signed(_T_904); // @[PositFMA.scala 60:76]
  assign _T_905 = $signed(sigA) * $signed(sigB); // @[PositFMA.scala 61:25]
  assign sigP = $unsigned(_T_905); // @[PositFMA.scala 61:33]
  assign head2 = sigP[51:50]; // @[PositFMA.scala 62:28]
  assign _T_906 = head2[1]; // @[PositFMA.scala 63:31]
  assign _T_907 = ~ _T_906; // @[PositFMA.scala 63:25]
  assign _T_908 = head2[0]; // @[PositFMA.scala 63:42]
  assign addTwo = _T_907 & _T_908; // @[PositFMA.scala 63:35]
  assign _T_909 = sigP[51]; // @[PositFMA.scala 65:23]
  assign _T_910 = sigP[49]; // @[PositFMA.scala 65:49]
  assign addOne = _T_909 ^ _T_910; // @[PositFMA.scala 65:43]
  assign _T_911 = {addTwo,addOne}; // @[Cat.scala 29:58]
  assign expBias = {1'b0,$signed(_T_911)}; // @[PositFMA.scala 66:39]
  assign mulSign = sigP[51:51]; // @[PositFMA.scala 67:28]
  assign _T_912 = $signed(decA_scale) + $signed(decB_scale); // @[PositFMA.scala 69:30]
  assign _GEN_12 = {{7{expBias[2]}},expBias}; // @[PositFMA.scala 69:44]
  assign _T_914 = $signed(_T_912) + $signed(_GEN_12); // @[PositFMA.scala 69:44]
  assign mulScale = $signed(_T_914); // @[PositFMA.scala 69:44]
  assign _T_915 = sigP[49:0]; // @[PositFMA.scala 72:29]
  assign _T_916 = sigP[48:0]; // @[PositFMA.scala 73:29]
  assign _T_917 = {_T_916, 1'h0}; // @[PositFMA.scala 73:48]
  assign mulSigTmp = addOne ? _T_915 : _T_917; // @[PositFMA.scala 70:22]
  assign _T_919 = mulSigTmp[49:49]; // @[PositFMA.scala 77:39]
  assign _T_920 = _T_919 | addTwo; // @[PositFMA.scala 77:43]
  assign _T_921 = mulSigTmp[48:0]; // @[PositFMA.scala 78:39]
  assign mulSig = {mulSign,_T_920,_T_921}; // @[Cat.scala 29:58]
  assign _T_947 = ~ addSign_phase2; // @[PositFMA.scala 107:29]
  assign _T_948 = ~ addZero_phase2; // @[PositFMA.scala 107:47]
  assign _T_949 = _T_947 & _T_948; // @[PositFMA.scala 107:45]
  assign extAddSig = {addSign_phase2,_T_949,addFrac_phase2,25'h0}; // @[Cat.scala 29:58]
  assign _GEN_13 = {{1{addScale_phase2[8]}},addScale_phase2}; // @[PositFMA.scala 111:39]
  assign mulGreater = $signed(mulScale_phase2) > $signed(_GEN_13); // @[PositFMA.scala 111:39]
  assign greaterScale = mulGreater ? $signed(mulScale_phase2) : $signed({{1{addScale_phase2[8]}},addScale_phase2}); // @[PositFMA.scala 112:26]
  assign smallerScale = mulGreater ? $signed({{1{addScale_phase2[8]}},addScale_phase2}) : $signed(mulScale_phase2); // @[PositFMA.scala 113:26]
  assign _T_953 = $signed(greaterScale) - $signed(smallerScale); // @[PositFMA.scala 114:36]
  assign scaleDiff = $signed(_T_953); // @[PositFMA.scala 114:36]
  assign greaterSig = mulGreater ? mulSig_phase2 : extAddSig; // @[PositFMA.scala 115:26]
  assign smallerSigTmp = mulGreater ? extAddSig : mulSig_phase2; // @[PositFMA.scala 116:26]
  assign _T_954 = $unsigned(scaleDiff); // @[PositFMA.scala 117:69]
  assign _T_955 = _T_954 < 10'h33; // @[Shift.scala 39:24]
  assign _T_956 = _T_954[5:0]; // @[Shift.scala 40:44]
  assign _T_957 = smallerSigTmp[50:32]; // @[Shift.scala 90:30]
  assign _T_958 = smallerSigTmp[31:0]; // @[Shift.scala 90:48]
  assign _T_959 = _T_958 != 32'h0; // @[Shift.scala 90:57]
  assign _GEN_14 = {{18'd0}, _T_959}; // @[Shift.scala 90:39]
  assign _T_960 = _T_957 | _GEN_14; // @[Shift.scala 90:39]
  assign _T_961 = _T_956[5]; // @[Shift.scala 12:21]
  assign _T_962 = smallerSigTmp[50]; // @[Shift.scala 12:21]
  assign _T_964 = _T_962 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 71:12]
  assign _T_965 = {_T_964,_T_960}; // @[Cat.scala 29:58]
  assign _T_966 = _T_961 ? _T_965 : smallerSigTmp; // @[Shift.scala 91:22]
  assign _T_967 = _T_956[4:0]; // @[Shift.scala 92:77]
  assign _T_968 = _T_966[50:16]; // @[Shift.scala 90:30]
  assign _T_969 = _T_966[15:0]; // @[Shift.scala 90:48]
  assign _T_970 = _T_969 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_15 = {{34'd0}, _T_970}; // @[Shift.scala 90:39]
  assign _T_971 = _T_968 | _GEN_15; // @[Shift.scala 90:39]
  assign _T_972 = _T_967[4]; // @[Shift.scala 12:21]
  assign _T_973 = _T_966[50]; // @[Shift.scala 12:21]
  assign _T_975 = _T_973 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_976 = {_T_975,_T_971}; // @[Cat.scala 29:58]
  assign _T_977 = _T_972 ? _T_976 : _T_966; // @[Shift.scala 91:22]
  assign _T_978 = _T_967[3:0]; // @[Shift.scala 92:77]
  assign _T_979 = _T_977[50:8]; // @[Shift.scala 90:30]
  assign _T_980 = _T_977[7:0]; // @[Shift.scala 90:48]
  assign _T_981 = _T_980 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_16 = {{42'd0}, _T_981}; // @[Shift.scala 90:39]
  assign _T_982 = _T_979 | _GEN_16; // @[Shift.scala 90:39]
  assign _T_983 = _T_978[3]; // @[Shift.scala 12:21]
  assign _T_984 = _T_977[50]; // @[Shift.scala 12:21]
  assign _T_986 = _T_984 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_987 = {_T_986,_T_982}; // @[Cat.scala 29:58]
  assign _T_988 = _T_983 ? _T_987 : _T_977; // @[Shift.scala 91:22]
  assign _T_989 = _T_978[2:0]; // @[Shift.scala 92:77]
  assign _T_990 = _T_988[50:4]; // @[Shift.scala 90:30]
  assign _T_991 = _T_988[3:0]; // @[Shift.scala 90:48]
  assign _T_992 = _T_991 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_17 = {{46'd0}, _T_992}; // @[Shift.scala 90:39]
  assign _T_993 = _T_990 | _GEN_17; // @[Shift.scala 90:39]
  assign _T_994 = _T_989[2]; // @[Shift.scala 12:21]
  assign _T_995 = _T_988[50]; // @[Shift.scala 12:21]
  assign _T_997 = _T_995 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_998 = {_T_997,_T_993}; // @[Cat.scala 29:58]
  assign _T_999 = _T_994 ? _T_998 : _T_988; // @[Shift.scala 91:22]
  assign _T_1000 = _T_989[1:0]; // @[Shift.scala 92:77]
  assign _T_1001 = _T_999[50:2]; // @[Shift.scala 90:30]
  assign _T_1002 = _T_999[1:0]; // @[Shift.scala 90:48]
  assign _T_1003 = _T_1002 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_18 = {{48'd0}, _T_1003}; // @[Shift.scala 90:39]
  assign _T_1004 = _T_1001 | _GEN_18; // @[Shift.scala 90:39]
  assign _T_1005 = _T_1000[1]; // @[Shift.scala 12:21]
  assign _T_1006 = _T_999[50]; // @[Shift.scala 12:21]
  assign _T_1008 = _T_1006 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_1009 = {_T_1008,_T_1004}; // @[Cat.scala 29:58]
  assign _T_1010 = _T_1005 ? _T_1009 : _T_999; // @[Shift.scala 91:22]
  assign _T_1011 = _T_1000[0:0]; // @[Shift.scala 92:77]
  assign _T_1012 = _T_1010[50:1]; // @[Shift.scala 90:30]
  assign _T_1013 = _T_1010[0:0]; // @[Shift.scala 90:48]
  assign _GEN_19 = {{49'd0}, _T_1013}; // @[Shift.scala 90:39]
  assign _T_1015 = _T_1012 | _GEN_19; // @[Shift.scala 90:39]
  assign _T_1017 = _T_1010[50]; // @[Shift.scala 12:21]
  assign _T_1018 = {_T_1017,_T_1015}; // @[Cat.scala 29:58]
  assign _T_1019 = _T_1011 ? _T_1018 : _T_1010; // @[Shift.scala 91:22]
  assign _T_1022 = _T_962 ? 51'h7ffffffffffff : 51'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_955 ? _T_1019 : _T_1022; // @[Shift.scala 39:10]
  assign rawSumSig = greaterSig + smallerSig; // @[PositFMA.scala 118:34]
  assign _T_1023 = mulSig_phase2[50:50]; // @[PositFMA.scala 119:42]
  assign _T_1024 = _T_1023 ^ addSign_phase2; // @[PositFMA.scala 119:46]
  assign _T_1025 = rawSumSig[51:51]; // @[PositFMA.scala 119:79]
  assign sumSign = _T_1024 ^ _T_1025; // @[PositFMA.scala 119:63]
  assign _T_1027 = greaterSig + smallerSig; // @[PositFMA.scala 120:50]
  assign signSumSig = {sumSign,_T_1027}; // @[Cat.scala 29:58]
  assign _T_1028 = signSumSig[51:1]; // @[PositFMA.scala 124:33]
  assign _T_1029 = signSumSig[50:0]; // @[PositFMA.scala 124:68]
  assign sumXor = _T_1028 ^ _T_1029; // @[PositFMA.scala 124:51]
  assign _T_1030 = sumXor[50:19]; // @[LZD.scala 43:32]
  assign _T_1031 = _T_1030[31:16]; // @[LZD.scala 43:32]
  assign _T_1032 = _T_1031[15:8]; // @[LZD.scala 43:32]
  assign _T_1033 = _T_1032[7:4]; // @[LZD.scala 43:32]
  assign _T_1034 = _T_1033[3:2]; // @[LZD.scala 43:32]
  assign _T_1035 = _T_1034 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1036 = _T_1034[1]; // @[LZD.scala 39:21]
  assign _T_1037 = _T_1034[0]; // @[LZD.scala 39:30]
  assign _T_1038 = ~ _T_1037; // @[LZD.scala 39:27]
  assign _T_1039 = _T_1036 | _T_1038; // @[LZD.scala 39:25]
  assign _T_1040 = {_T_1035,_T_1039}; // @[Cat.scala 29:58]
  assign _T_1041 = _T_1033[1:0]; // @[LZD.scala 44:32]
  assign _T_1042 = _T_1041 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1043 = _T_1041[1]; // @[LZD.scala 39:21]
  assign _T_1044 = _T_1041[0]; // @[LZD.scala 39:30]
  assign _T_1045 = ~ _T_1044; // @[LZD.scala 39:27]
  assign _T_1046 = _T_1043 | _T_1045; // @[LZD.scala 39:25]
  assign _T_1047 = {_T_1042,_T_1046}; // @[Cat.scala 29:58]
  assign _T_1048 = _T_1040[1]; // @[Shift.scala 12:21]
  assign _T_1049 = _T_1047[1]; // @[Shift.scala 12:21]
  assign _T_1050 = _T_1048 | _T_1049; // @[LZD.scala 49:16]
  assign _T_1051 = ~ _T_1049; // @[LZD.scala 49:27]
  assign _T_1052 = _T_1048 | _T_1051; // @[LZD.scala 49:25]
  assign _T_1053 = _T_1040[0:0]; // @[LZD.scala 49:47]
  assign _T_1054 = _T_1047[0:0]; // @[LZD.scala 49:59]
  assign _T_1055 = _T_1048 ? _T_1053 : _T_1054; // @[LZD.scala 49:35]
  assign _T_1057 = {_T_1050,_T_1052,_T_1055}; // @[Cat.scala 29:58]
  assign _T_1058 = _T_1032[3:0]; // @[LZD.scala 44:32]
  assign _T_1059 = _T_1058[3:2]; // @[LZD.scala 43:32]
  assign _T_1060 = _T_1059 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1061 = _T_1059[1]; // @[LZD.scala 39:21]
  assign _T_1062 = _T_1059[0]; // @[LZD.scala 39:30]
  assign _T_1063 = ~ _T_1062; // @[LZD.scala 39:27]
  assign _T_1064 = _T_1061 | _T_1063; // @[LZD.scala 39:25]
  assign _T_1065 = {_T_1060,_T_1064}; // @[Cat.scala 29:58]
  assign _T_1066 = _T_1058[1:0]; // @[LZD.scala 44:32]
  assign _T_1067 = _T_1066 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1068 = _T_1066[1]; // @[LZD.scala 39:21]
  assign _T_1069 = _T_1066[0]; // @[LZD.scala 39:30]
  assign _T_1070 = ~ _T_1069; // @[LZD.scala 39:27]
  assign _T_1071 = _T_1068 | _T_1070; // @[LZD.scala 39:25]
  assign _T_1072 = {_T_1067,_T_1071}; // @[Cat.scala 29:58]
  assign _T_1073 = _T_1065[1]; // @[Shift.scala 12:21]
  assign _T_1074 = _T_1072[1]; // @[Shift.scala 12:21]
  assign _T_1075 = _T_1073 | _T_1074; // @[LZD.scala 49:16]
  assign _T_1076 = ~ _T_1074; // @[LZD.scala 49:27]
  assign _T_1077 = _T_1073 | _T_1076; // @[LZD.scala 49:25]
  assign _T_1078 = _T_1065[0:0]; // @[LZD.scala 49:47]
  assign _T_1079 = _T_1072[0:0]; // @[LZD.scala 49:59]
  assign _T_1080 = _T_1073 ? _T_1078 : _T_1079; // @[LZD.scala 49:35]
  assign _T_1082 = {_T_1075,_T_1077,_T_1080}; // @[Cat.scala 29:58]
  assign _T_1083 = _T_1057[2]; // @[Shift.scala 12:21]
  assign _T_1084 = _T_1082[2]; // @[Shift.scala 12:21]
  assign _T_1085 = _T_1083 | _T_1084; // @[LZD.scala 49:16]
  assign _T_1086 = ~ _T_1084; // @[LZD.scala 49:27]
  assign _T_1087 = _T_1083 | _T_1086; // @[LZD.scala 49:25]
  assign _T_1088 = _T_1057[1:0]; // @[LZD.scala 49:47]
  assign _T_1089 = _T_1082[1:0]; // @[LZD.scala 49:59]
  assign _T_1090 = _T_1083 ? _T_1088 : _T_1089; // @[LZD.scala 49:35]
  assign _T_1092 = {_T_1085,_T_1087,_T_1090}; // @[Cat.scala 29:58]
  assign _T_1093 = _T_1031[7:0]; // @[LZD.scala 44:32]
  assign _T_1094 = _T_1093[7:4]; // @[LZD.scala 43:32]
  assign _T_1095 = _T_1094[3:2]; // @[LZD.scala 43:32]
  assign _T_1096 = _T_1095 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1097 = _T_1095[1]; // @[LZD.scala 39:21]
  assign _T_1098 = _T_1095[0]; // @[LZD.scala 39:30]
  assign _T_1099 = ~ _T_1098; // @[LZD.scala 39:27]
  assign _T_1100 = _T_1097 | _T_1099; // @[LZD.scala 39:25]
  assign _T_1101 = {_T_1096,_T_1100}; // @[Cat.scala 29:58]
  assign _T_1102 = _T_1094[1:0]; // @[LZD.scala 44:32]
  assign _T_1103 = _T_1102 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1104 = _T_1102[1]; // @[LZD.scala 39:21]
  assign _T_1105 = _T_1102[0]; // @[LZD.scala 39:30]
  assign _T_1106 = ~ _T_1105; // @[LZD.scala 39:27]
  assign _T_1107 = _T_1104 | _T_1106; // @[LZD.scala 39:25]
  assign _T_1108 = {_T_1103,_T_1107}; // @[Cat.scala 29:58]
  assign _T_1109 = _T_1101[1]; // @[Shift.scala 12:21]
  assign _T_1110 = _T_1108[1]; // @[Shift.scala 12:21]
  assign _T_1111 = _T_1109 | _T_1110; // @[LZD.scala 49:16]
  assign _T_1112 = ~ _T_1110; // @[LZD.scala 49:27]
  assign _T_1113 = _T_1109 | _T_1112; // @[LZD.scala 49:25]
  assign _T_1114 = _T_1101[0:0]; // @[LZD.scala 49:47]
  assign _T_1115 = _T_1108[0:0]; // @[LZD.scala 49:59]
  assign _T_1116 = _T_1109 ? _T_1114 : _T_1115; // @[LZD.scala 49:35]
  assign _T_1118 = {_T_1111,_T_1113,_T_1116}; // @[Cat.scala 29:58]
  assign _T_1119 = _T_1093[3:0]; // @[LZD.scala 44:32]
  assign _T_1120 = _T_1119[3:2]; // @[LZD.scala 43:32]
  assign _T_1121 = _T_1120 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1122 = _T_1120[1]; // @[LZD.scala 39:21]
  assign _T_1123 = _T_1120[0]; // @[LZD.scala 39:30]
  assign _T_1124 = ~ _T_1123; // @[LZD.scala 39:27]
  assign _T_1125 = _T_1122 | _T_1124; // @[LZD.scala 39:25]
  assign _T_1126 = {_T_1121,_T_1125}; // @[Cat.scala 29:58]
  assign _T_1127 = _T_1119[1:0]; // @[LZD.scala 44:32]
  assign _T_1128 = _T_1127 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1129 = _T_1127[1]; // @[LZD.scala 39:21]
  assign _T_1130 = _T_1127[0]; // @[LZD.scala 39:30]
  assign _T_1131 = ~ _T_1130; // @[LZD.scala 39:27]
  assign _T_1132 = _T_1129 | _T_1131; // @[LZD.scala 39:25]
  assign _T_1133 = {_T_1128,_T_1132}; // @[Cat.scala 29:58]
  assign _T_1134 = _T_1126[1]; // @[Shift.scala 12:21]
  assign _T_1135 = _T_1133[1]; // @[Shift.scala 12:21]
  assign _T_1136 = _T_1134 | _T_1135; // @[LZD.scala 49:16]
  assign _T_1137 = ~ _T_1135; // @[LZD.scala 49:27]
  assign _T_1138 = _T_1134 | _T_1137; // @[LZD.scala 49:25]
  assign _T_1139 = _T_1126[0:0]; // @[LZD.scala 49:47]
  assign _T_1140 = _T_1133[0:0]; // @[LZD.scala 49:59]
  assign _T_1141 = _T_1134 ? _T_1139 : _T_1140; // @[LZD.scala 49:35]
  assign _T_1143 = {_T_1136,_T_1138,_T_1141}; // @[Cat.scala 29:58]
  assign _T_1144 = _T_1118[2]; // @[Shift.scala 12:21]
  assign _T_1145 = _T_1143[2]; // @[Shift.scala 12:21]
  assign _T_1146 = _T_1144 | _T_1145; // @[LZD.scala 49:16]
  assign _T_1147 = ~ _T_1145; // @[LZD.scala 49:27]
  assign _T_1148 = _T_1144 | _T_1147; // @[LZD.scala 49:25]
  assign _T_1149 = _T_1118[1:0]; // @[LZD.scala 49:47]
  assign _T_1150 = _T_1143[1:0]; // @[LZD.scala 49:59]
  assign _T_1151 = _T_1144 ? _T_1149 : _T_1150; // @[LZD.scala 49:35]
  assign _T_1153 = {_T_1146,_T_1148,_T_1151}; // @[Cat.scala 29:58]
  assign _T_1154 = _T_1092[3]; // @[Shift.scala 12:21]
  assign _T_1155 = _T_1153[3]; // @[Shift.scala 12:21]
  assign _T_1156 = _T_1154 | _T_1155; // @[LZD.scala 49:16]
  assign _T_1157 = ~ _T_1155; // @[LZD.scala 49:27]
  assign _T_1158 = _T_1154 | _T_1157; // @[LZD.scala 49:25]
  assign _T_1159 = _T_1092[2:0]; // @[LZD.scala 49:47]
  assign _T_1160 = _T_1153[2:0]; // @[LZD.scala 49:59]
  assign _T_1161 = _T_1154 ? _T_1159 : _T_1160; // @[LZD.scala 49:35]
  assign _T_1163 = {_T_1156,_T_1158,_T_1161}; // @[Cat.scala 29:58]
  assign _T_1164 = _T_1030[15:0]; // @[LZD.scala 44:32]
  assign _T_1165 = _T_1164[15:8]; // @[LZD.scala 43:32]
  assign _T_1166 = _T_1165[7:4]; // @[LZD.scala 43:32]
  assign _T_1167 = _T_1166[3:2]; // @[LZD.scala 43:32]
  assign _T_1168 = _T_1167 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1169 = _T_1167[1]; // @[LZD.scala 39:21]
  assign _T_1170 = _T_1167[0]; // @[LZD.scala 39:30]
  assign _T_1171 = ~ _T_1170; // @[LZD.scala 39:27]
  assign _T_1172 = _T_1169 | _T_1171; // @[LZD.scala 39:25]
  assign _T_1173 = {_T_1168,_T_1172}; // @[Cat.scala 29:58]
  assign _T_1174 = _T_1166[1:0]; // @[LZD.scala 44:32]
  assign _T_1175 = _T_1174 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1176 = _T_1174[1]; // @[LZD.scala 39:21]
  assign _T_1177 = _T_1174[0]; // @[LZD.scala 39:30]
  assign _T_1178 = ~ _T_1177; // @[LZD.scala 39:27]
  assign _T_1179 = _T_1176 | _T_1178; // @[LZD.scala 39:25]
  assign _T_1180 = {_T_1175,_T_1179}; // @[Cat.scala 29:58]
  assign _T_1181 = _T_1173[1]; // @[Shift.scala 12:21]
  assign _T_1182 = _T_1180[1]; // @[Shift.scala 12:21]
  assign _T_1183 = _T_1181 | _T_1182; // @[LZD.scala 49:16]
  assign _T_1184 = ~ _T_1182; // @[LZD.scala 49:27]
  assign _T_1185 = _T_1181 | _T_1184; // @[LZD.scala 49:25]
  assign _T_1186 = _T_1173[0:0]; // @[LZD.scala 49:47]
  assign _T_1187 = _T_1180[0:0]; // @[LZD.scala 49:59]
  assign _T_1188 = _T_1181 ? _T_1186 : _T_1187; // @[LZD.scala 49:35]
  assign _T_1190 = {_T_1183,_T_1185,_T_1188}; // @[Cat.scala 29:58]
  assign _T_1191 = _T_1165[3:0]; // @[LZD.scala 44:32]
  assign _T_1192 = _T_1191[3:2]; // @[LZD.scala 43:32]
  assign _T_1193 = _T_1192 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1194 = _T_1192[1]; // @[LZD.scala 39:21]
  assign _T_1195 = _T_1192[0]; // @[LZD.scala 39:30]
  assign _T_1196 = ~ _T_1195; // @[LZD.scala 39:27]
  assign _T_1197 = _T_1194 | _T_1196; // @[LZD.scala 39:25]
  assign _T_1198 = {_T_1193,_T_1197}; // @[Cat.scala 29:58]
  assign _T_1199 = _T_1191[1:0]; // @[LZD.scala 44:32]
  assign _T_1200 = _T_1199 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1201 = _T_1199[1]; // @[LZD.scala 39:21]
  assign _T_1202 = _T_1199[0]; // @[LZD.scala 39:30]
  assign _T_1203 = ~ _T_1202; // @[LZD.scala 39:27]
  assign _T_1204 = _T_1201 | _T_1203; // @[LZD.scala 39:25]
  assign _T_1205 = {_T_1200,_T_1204}; // @[Cat.scala 29:58]
  assign _T_1206 = _T_1198[1]; // @[Shift.scala 12:21]
  assign _T_1207 = _T_1205[1]; // @[Shift.scala 12:21]
  assign _T_1208 = _T_1206 | _T_1207; // @[LZD.scala 49:16]
  assign _T_1209 = ~ _T_1207; // @[LZD.scala 49:27]
  assign _T_1210 = _T_1206 | _T_1209; // @[LZD.scala 49:25]
  assign _T_1211 = _T_1198[0:0]; // @[LZD.scala 49:47]
  assign _T_1212 = _T_1205[0:0]; // @[LZD.scala 49:59]
  assign _T_1213 = _T_1206 ? _T_1211 : _T_1212; // @[LZD.scala 49:35]
  assign _T_1215 = {_T_1208,_T_1210,_T_1213}; // @[Cat.scala 29:58]
  assign _T_1216 = _T_1190[2]; // @[Shift.scala 12:21]
  assign _T_1217 = _T_1215[2]; // @[Shift.scala 12:21]
  assign _T_1218 = _T_1216 | _T_1217; // @[LZD.scala 49:16]
  assign _T_1219 = ~ _T_1217; // @[LZD.scala 49:27]
  assign _T_1220 = _T_1216 | _T_1219; // @[LZD.scala 49:25]
  assign _T_1221 = _T_1190[1:0]; // @[LZD.scala 49:47]
  assign _T_1222 = _T_1215[1:0]; // @[LZD.scala 49:59]
  assign _T_1223 = _T_1216 ? _T_1221 : _T_1222; // @[LZD.scala 49:35]
  assign _T_1225 = {_T_1218,_T_1220,_T_1223}; // @[Cat.scala 29:58]
  assign _T_1226 = _T_1164[7:0]; // @[LZD.scala 44:32]
  assign _T_1227 = _T_1226[7:4]; // @[LZD.scala 43:32]
  assign _T_1228 = _T_1227[3:2]; // @[LZD.scala 43:32]
  assign _T_1229 = _T_1228 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1230 = _T_1228[1]; // @[LZD.scala 39:21]
  assign _T_1231 = _T_1228[0]; // @[LZD.scala 39:30]
  assign _T_1232 = ~ _T_1231; // @[LZD.scala 39:27]
  assign _T_1233 = _T_1230 | _T_1232; // @[LZD.scala 39:25]
  assign _T_1234 = {_T_1229,_T_1233}; // @[Cat.scala 29:58]
  assign _T_1235 = _T_1227[1:0]; // @[LZD.scala 44:32]
  assign _T_1236 = _T_1235 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1237 = _T_1235[1]; // @[LZD.scala 39:21]
  assign _T_1238 = _T_1235[0]; // @[LZD.scala 39:30]
  assign _T_1239 = ~ _T_1238; // @[LZD.scala 39:27]
  assign _T_1240 = _T_1237 | _T_1239; // @[LZD.scala 39:25]
  assign _T_1241 = {_T_1236,_T_1240}; // @[Cat.scala 29:58]
  assign _T_1242 = _T_1234[1]; // @[Shift.scala 12:21]
  assign _T_1243 = _T_1241[1]; // @[Shift.scala 12:21]
  assign _T_1244 = _T_1242 | _T_1243; // @[LZD.scala 49:16]
  assign _T_1245 = ~ _T_1243; // @[LZD.scala 49:27]
  assign _T_1246 = _T_1242 | _T_1245; // @[LZD.scala 49:25]
  assign _T_1247 = _T_1234[0:0]; // @[LZD.scala 49:47]
  assign _T_1248 = _T_1241[0:0]; // @[LZD.scala 49:59]
  assign _T_1249 = _T_1242 ? _T_1247 : _T_1248; // @[LZD.scala 49:35]
  assign _T_1251 = {_T_1244,_T_1246,_T_1249}; // @[Cat.scala 29:58]
  assign _T_1252 = _T_1226[3:0]; // @[LZD.scala 44:32]
  assign _T_1253 = _T_1252[3:2]; // @[LZD.scala 43:32]
  assign _T_1254 = _T_1253 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1255 = _T_1253[1]; // @[LZD.scala 39:21]
  assign _T_1256 = _T_1253[0]; // @[LZD.scala 39:30]
  assign _T_1257 = ~ _T_1256; // @[LZD.scala 39:27]
  assign _T_1258 = _T_1255 | _T_1257; // @[LZD.scala 39:25]
  assign _T_1259 = {_T_1254,_T_1258}; // @[Cat.scala 29:58]
  assign _T_1260 = _T_1252[1:0]; // @[LZD.scala 44:32]
  assign _T_1261 = _T_1260 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1262 = _T_1260[1]; // @[LZD.scala 39:21]
  assign _T_1263 = _T_1260[0]; // @[LZD.scala 39:30]
  assign _T_1264 = ~ _T_1263; // @[LZD.scala 39:27]
  assign _T_1265 = _T_1262 | _T_1264; // @[LZD.scala 39:25]
  assign _T_1266 = {_T_1261,_T_1265}; // @[Cat.scala 29:58]
  assign _T_1267 = _T_1259[1]; // @[Shift.scala 12:21]
  assign _T_1268 = _T_1266[1]; // @[Shift.scala 12:21]
  assign _T_1269 = _T_1267 | _T_1268; // @[LZD.scala 49:16]
  assign _T_1270 = ~ _T_1268; // @[LZD.scala 49:27]
  assign _T_1271 = _T_1267 | _T_1270; // @[LZD.scala 49:25]
  assign _T_1272 = _T_1259[0:0]; // @[LZD.scala 49:47]
  assign _T_1273 = _T_1266[0:0]; // @[LZD.scala 49:59]
  assign _T_1274 = _T_1267 ? _T_1272 : _T_1273; // @[LZD.scala 49:35]
  assign _T_1276 = {_T_1269,_T_1271,_T_1274}; // @[Cat.scala 29:58]
  assign _T_1277 = _T_1251[2]; // @[Shift.scala 12:21]
  assign _T_1278 = _T_1276[2]; // @[Shift.scala 12:21]
  assign _T_1279 = _T_1277 | _T_1278; // @[LZD.scala 49:16]
  assign _T_1280 = ~ _T_1278; // @[LZD.scala 49:27]
  assign _T_1281 = _T_1277 | _T_1280; // @[LZD.scala 49:25]
  assign _T_1282 = _T_1251[1:0]; // @[LZD.scala 49:47]
  assign _T_1283 = _T_1276[1:0]; // @[LZD.scala 49:59]
  assign _T_1284 = _T_1277 ? _T_1282 : _T_1283; // @[LZD.scala 49:35]
  assign _T_1286 = {_T_1279,_T_1281,_T_1284}; // @[Cat.scala 29:58]
  assign _T_1287 = _T_1225[3]; // @[Shift.scala 12:21]
  assign _T_1288 = _T_1286[3]; // @[Shift.scala 12:21]
  assign _T_1289 = _T_1287 | _T_1288; // @[LZD.scala 49:16]
  assign _T_1290 = ~ _T_1288; // @[LZD.scala 49:27]
  assign _T_1291 = _T_1287 | _T_1290; // @[LZD.scala 49:25]
  assign _T_1292 = _T_1225[2:0]; // @[LZD.scala 49:47]
  assign _T_1293 = _T_1286[2:0]; // @[LZD.scala 49:59]
  assign _T_1294 = _T_1287 ? _T_1292 : _T_1293; // @[LZD.scala 49:35]
  assign _T_1296 = {_T_1289,_T_1291,_T_1294}; // @[Cat.scala 29:58]
  assign _T_1297 = _T_1163[4]; // @[Shift.scala 12:21]
  assign _T_1298 = _T_1296[4]; // @[Shift.scala 12:21]
  assign _T_1299 = _T_1297 | _T_1298; // @[LZD.scala 49:16]
  assign _T_1300 = ~ _T_1298; // @[LZD.scala 49:27]
  assign _T_1301 = _T_1297 | _T_1300; // @[LZD.scala 49:25]
  assign _T_1302 = _T_1163[3:0]; // @[LZD.scala 49:47]
  assign _T_1303 = _T_1296[3:0]; // @[LZD.scala 49:59]
  assign _T_1304 = _T_1297 ? _T_1302 : _T_1303; // @[LZD.scala 49:35]
  assign _T_1306 = {_T_1299,_T_1301,_T_1304}; // @[Cat.scala 29:58]
  assign _T_1307 = sumXor[18:0]; // @[LZD.scala 44:32]
  assign _T_1308 = _T_1307[18:3]; // @[LZD.scala 43:32]
  assign _T_1309 = _T_1308[15:8]; // @[LZD.scala 43:32]
  assign _T_1310 = _T_1309[7:4]; // @[LZD.scala 43:32]
  assign _T_1311 = _T_1310[3:2]; // @[LZD.scala 43:32]
  assign _T_1312 = _T_1311 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1313 = _T_1311[1]; // @[LZD.scala 39:21]
  assign _T_1314 = _T_1311[0]; // @[LZD.scala 39:30]
  assign _T_1315 = ~ _T_1314; // @[LZD.scala 39:27]
  assign _T_1316 = _T_1313 | _T_1315; // @[LZD.scala 39:25]
  assign _T_1317 = {_T_1312,_T_1316}; // @[Cat.scala 29:58]
  assign _T_1318 = _T_1310[1:0]; // @[LZD.scala 44:32]
  assign _T_1319 = _T_1318 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1320 = _T_1318[1]; // @[LZD.scala 39:21]
  assign _T_1321 = _T_1318[0]; // @[LZD.scala 39:30]
  assign _T_1322 = ~ _T_1321; // @[LZD.scala 39:27]
  assign _T_1323 = _T_1320 | _T_1322; // @[LZD.scala 39:25]
  assign _T_1324 = {_T_1319,_T_1323}; // @[Cat.scala 29:58]
  assign _T_1325 = _T_1317[1]; // @[Shift.scala 12:21]
  assign _T_1326 = _T_1324[1]; // @[Shift.scala 12:21]
  assign _T_1327 = _T_1325 | _T_1326; // @[LZD.scala 49:16]
  assign _T_1328 = ~ _T_1326; // @[LZD.scala 49:27]
  assign _T_1329 = _T_1325 | _T_1328; // @[LZD.scala 49:25]
  assign _T_1330 = _T_1317[0:0]; // @[LZD.scala 49:47]
  assign _T_1331 = _T_1324[0:0]; // @[LZD.scala 49:59]
  assign _T_1332 = _T_1325 ? _T_1330 : _T_1331; // @[LZD.scala 49:35]
  assign _T_1334 = {_T_1327,_T_1329,_T_1332}; // @[Cat.scala 29:58]
  assign _T_1335 = _T_1309[3:0]; // @[LZD.scala 44:32]
  assign _T_1336 = _T_1335[3:2]; // @[LZD.scala 43:32]
  assign _T_1337 = _T_1336 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1338 = _T_1336[1]; // @[LZD.scala 39:21]
  assign _T_1339 = _T_1336[0]; // @[LZD.scala 39:30]
  assign _T_1340 = ~ _T_1339; // @[LZD.scala 39:27]
  assign _T_1341 = _T_1338 | _T_1340; // @[LZD.scala 39:25]
  assign _T_1342 = {_T_1337,_T_1341}; // @[Cat.scala 29:58]
  assign _T_1343 = _T_1335[1:0]; // @[LZD.scala 44:32]
  assign _T_1344 = _T_1343 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1345 = _T_1343[1]; // @[LZD.scala 39:21]
  assign _T_1346 = _T_1343[0]; // @[LZD.scala 39:30]
  assign _T_1347 = ~ _T_1346; // @[LZD.scala 39:27]
  assign _T_1348 = _T_1345 | _T_1347; // @[LZD.scala 39:25]
  assign _T_1349 = {_T_1344,_T_1348}; // @[Cat.scala 29:58]
  assign _T_1350 = _T_1342[1]; // @[Shift.scala 12:21]
  assign _T_1351 = _T_1349[1]; // @[Shift.scala 12:21]
  assign _T_1352 = _T_1350 | _T_1351; // @[LZD.scala 49:16]
  assign _T_1353 = ~ _T_1351; // @[LZD.scala 49:27]
  assign _T_1354 = _T_1350 | _T_1353; // @[LZD.scala 49:25]
  assign _T_1355 = _T_1342[0:0]; // @[LZD.scala 49:47]
  assign _T_1356 = _T_1349[0:0]; // @[LZD.scala 49:59]
  assign _T_1357 = _T_1350 ? _T_1355 : _T_1356; // @[LZD.scala 49:35]
  assign _T_1359 = {_T_1352,_T_1354,_T_1357}; // @[Cat.scala 29:58]
  assign _T_1360 = _T_1334[2]; // @[Shift.scala 12:21]
  assign _T_1361 = _T_1359[2]; // @[Shift.scala 12:21]
  assign _T_1362 = _T_1360 | _T_1361; // @[LZD.scala 49:16]
  assign _T_1363 = ~ _T_1361; // @[LZD.scala 49:27]
  assign _T_1364 = _T_1360 | _T_1363; // @[LZD.scala 49:25]
  assign _T_1365 = _T_1334[1:0]; // @[LZD.scala 49:47]
  assign _T_1366 = _T_1359[1:0]; // @[LZD.scala 49:59]
  assign _T_1367 = _T_1360 ? _T_1365 : _T_1366; // @[LZD.scala 49:35]
  assign _T_1369 = {_T_1362,_T_1364,_T_1367}; // @[Cat.scala 29:58]
  assign _T_1370 = _T_1308[7:0]; // @[LZD.scala 44:32]
  assign _T_1371 = _T_1370[7:4]; // @[LZD.scala 43:32]
  assign _T_1372 = _T_1371[3:2]; // @[LZD.scala 43:32]
  assign _T_1373 = _T_1372 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1374 = _T_1372[1]; // @[LZD.scala 39:21]
  assign _T_1375 = _T_1372[0]; // @[LZD.scala 39:30]
  assign _T_1376 = ~ _T_1375; // @[LZD.scala 39:27]
  assign _T_1377 = _T_1374 | _T_1376; // @[LZD.scala 39:25]
  assign _T_1378 = {_T_1373,_T_1377}; // @[Cat.scala 29:58]
  assign _T_1379 = _T_1371[1:0]; // @[LZD.scala 44:32]
  assign _T_1380 = _T_1379 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1381 = _T_1379[1]; // @[LZD.scala 39:21]
  assign _T_1382 = _T_1379[0]; // @[LZD.scala 39:30]
  assign _T_1383 = ~ _T_1382; // @[LZD.scala 39:27]
  assign _T_1384 = _T_1381 | _T_1383; // @[LZD.scala 39:25]
  assign _T_1385 = {_T_1380,_T_1384}; // @[Cat.scala 29:58]
  assign _T_1386 = _T_1378[1]; // @[Shift.scala 12:21]
  assign _T_1387 = _T_1385[1]; // @[Shift.scala 12:21]
  assign _T_1388 = _T_1386 | _T_1387; // @[LZD.scala 49:16]
  assign _T_1389 = ~ _T_1387; // @[LZD.scala 49:27]
  assign _T_1390 = _T_1386 | _T_1389; // @[LZD.scala 49:25]
  assign _T_1391 = _T_1378[0:0]; // @[LZD.scala 49:47]
  assign _T_1392 = _T_1385[0:0]; // @[LZD.scala 49:59]
  assign _T_1393 = _T_1386 ? _T_1391 : _T_1392; // @[LZD.scala 49:35]
  assign _T_1395 = {_T_1388,_T_1390,_T_1393}; // @[Cat.scala 29:58]
  assign _T_1396 = _T_1370[3:0]; // @[LZD.scala 44:32]
  assign _T_1397 = _T_1396[3:2]; // @[LZD.scala 43:32]
  assign _T_1398 = _T_1397 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1399 = _T_1397[1]; // @[LZD.scala 39:21]
  assign _T_1400 = _T_1397[0]; // @[LZD.scala 39:30]
  assign _T_1401 = ~ _T_1400; // @[LZD.scala 39:27]
  assign _T_1402 = _T_1399 | _T_1401; // @[LZD.scala 39:25]
  assign _T_1403 = {_T_1398,_T_1402}; // @[Cat.scala 29:58]
  assign _T_1404 = _T_1396[1:0]; // @[LZD.scala 44:32]
  assign _T_1405 = _T_1404 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1406 = _T_1404[1]; // @[LZD.scala 39:21]
  assign _T_1407 = _T_1404[0]; // @[LZD.scala 39:30]
  assign _T_1408 = ~ _T_1407; // @[LZD.scala 39:27]
  assign _T_1409 = _T_1406 | _T_1408; // @[LZD.scala 39:25]
  assign _T_1410 = {_T_1405,_T_1409}; // @[Cat.scala 29:58]
  assign _T_1411 = _T_1403[1]; // @[Shift.scala 12:21]
  assign _T_1412 = _T_1410[1]; // @[Shift.scala 12:21]
  assign _T_1413 = _T_1411 | _T_1412; // @[LZD.scala 49:16]
  assign _T_1414 = ~ _T_1412; // @[LZD.scala 49:27]
  assign _T_1415 = _T_1411 | _T_1414; // @[LZD.scala 49:25]
  assign _T_1416 = _T_1403[0:0]; // @[LZD.scala 49:47]
  assign _T_1417 = _T_1410[0:0]; // @[LZD.scala 49:59]
  assign _T_1418 = _T_1411 ? _T_1416 : _T_1417; // @[LZD.scala 49:35]
  assign _T_1420 = {_T_1413,_T_1415,_T_1418}; // @[Cat.scala 29:58]
  assign _T_1421 = _T_1395[2]; // @[Shift.scala 12:21]
  assign _T_1422 = _T_1420[2]; // @[Shift.scala 12:21]
  assign _T_1423 = _T_1421 | _T_1422; // @[LZD.scala 49:16]
  assign _T_1424 = ~ _T_1422; // @[LZD.scala 49:27]
  assign _T_1425 = _T_1421 | _T_1424; // @[LZD.scala 49:25]
  assign _T_1426 = _T_1395[1:0]; // @[LZD.scala 49:47]
  assign _T_1427 = _T_1420[1:0]; // @[LZD.scala 49:59]
  assign _T_1428 = _T_1421 ? _T_1426 : _T_1427; // @[LZD.scala 49:35]
  assign _T_1430 = {_T_1423,_T_1425,_T_1428}; // @[Cat.scala 29:58]
  assign _T_1431 = _T_1369[3]; // @[Shift.scala 12:21]
  assign _T_1432 = _T_1430[3]; // @[Shift.scala 12:21]
  assign _T_1433 = _T_1431 | _T_1432; // @[LZD.scala 49:16]
  assign _T_1434 = ~ _T_1432; // @[LZD.scala 49:27]
  assign _T_1435 = _T_1431 | _T_1434; // @[LZD.scala 49:25]
  assign _T_1436 = _T_1369[2:0]; // @[LZD.scala 49:47]
  assign _T_1437 = _T_1430[2:0]; // @[LZD.scala 49:59]
  assign _T_1438 = _T_1431 ? _T_1436 : _T_1437; // @[LZD.scala 49:35]
  assign _T_1440 = {_T_1433,_T_1435,_T_1438}; // @[Cat.scala 29:58]
  assign _T_1441 = _T_1307[2:0]; // @[LZD.scala 44:32]
  assign _T_1442 = _T_1441[2:1]; // @[LZD.scala 43:32]
  assign _T_1443 = _T_1442 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1444 = _T_1442[1]; // @[LZD.scala 39:21]
  assign _T_1445 = _T_1442[0]; // @[LZD.scala 39:30]
  assign _T_1446 = ~ _T_1445; // @[LZD.scala 39:27]
  assign _T_1447 = _T_1444 | _T_1446; // @[LZD.scala 39:25]
  assign _T_1448 = {_T_1443,_T_1447}; // @[Cat.scala 29:58]
  assign _T_1449 = _T_1441[0:0]; // @[LZD.scala 44:32]
  assign _T_1451 = _T_1448[1]; // @[Shift.scala 12:21]
  assign _T_1453 = _T_1448[0:0]; // @[LZD.scala 55:32]
  assign _T_1454 = _T_1451 ? _T_1453 : _T_1449; // @[LZD.scala 55:20]
  assign _T_1456 = _T_1440[4]; // @[Shift.scala 12:21]
  assign _T_1459 = {2'h3,_T_1451,_T_1454}; // @[Cat.scala 29:58]
  assign _T_1460 = _T_1440[3:0]; // @[LZD.scala 55:32]
  assign _T_1461 = _T_1456 ? _T_1460 : _T_1459; // @[LZD.scala 55:20]
  assign _T_1462 = {_T_1456,_T_1461}; // @[Cat.scala 29:58]
  assign _T_1463 = _T_1306[5]; // @[Shift.scala 12:21]
  assign _T_1465 = _T_1306[4:0]; // @[LZD.scala 55:32]
  assign _T_1466 = _T_1463 ? _T_1465 : _T_1462; // @[LZD.scala 55:20]
  assign sumLZD = {_T_1463,_T_1466}; // @[Cat.scala 29:58]
  assign shiftValue = ~ sumLZD; // @[PositFMA.scala 126:24]
  assign _T_1467 = signSumSig[49:0]; // @[PositFMA.scala 127:38]
  assign _T_1468 = shiftValue < 6'h32; // @[Shift.scala 16:24]
  assign _T_1470 = shiftValue[5]; // @[Shift.scala 12:21]
  assign _T_1471 = _T_1467[17:0]; // @[Shift.scala 64:52]
  assign _T_1473 = {_T_1471,32'h0}; // @[Cat.scala 29:58]
  assign _T_1474 = _T_1470 ? _T_1473 : _T_1467; // @[Shift.scala 64:27]
  assign _T_1475 = shiftValue[4:0]; // @[Shift.scala 66:70]
  assign _T_1476 = _T_1475[4]; // @[Shift.scala 12:21]
  assign _T_1477 = _T_1474[33:0]; // @[Shift.scala 64:52]
  assign _T_1479 = {_T_1477,16'h0}; // @[Cat.scala 29:58]
  assign _T_1480 = _T_1476 ? _T_1479 : _T_1474; // @[Shift.scala 64:27]
  assign _T_1481 = _T_1475[3:0]; // @[Shift.scala 66:70]
  assign _T_1482 = _T_1481[3]; // @[Shift.scala 12:21]
  assign _T_1483 = _T_1480[41:0]; // @[Shift.scala 64:52]
  assign _T_1485 = {_T_1483,8'h0}; // @[Cat.scala 29:58]
  assign _T_1486 = _T_1482 ? _T_1485 : _T_1480; // @[Shift.scala 64:27]
  assign _T_1487 = _T_1481[2:0]; // @[Shift.scala 66:70]
  assign _T_1488 = _T_1487[2]; // @[Shift.scala 12:21]
  assign _T_1489 = _T_1486[45:0]; // @[Shift.scala 64:52]
  assign _T_1491 = {_T_1489,4'h0}; // @[Cat.scala 29:58]
  assign _T_1492 = _T_1488 ? _T_1491 : _T_1486; // @[Shift.scala 64:27]
  assign _T_1493 = _T_1487[1:0]; // @[Shift.scala 66:70]
  assign _T_1494 = _T_1493[1]; // @[Shift.scala 12:21]
  assign _T_1495 = _T_1492[47:0]; // @[Shift.scala 64:52]
  assign _T_1497 = {_T_1495,2'h0}; // @[Cat.scala 29:58]
  assign _T_1498 = _T_1494 ? _T_1497 : _T_1492; // @[Shift.scala 64:27]
  assign _T_1499 = _T_1493[0:0]; // @[Shift.scala 66:70]
  assign _T_1501 = _T_1498[48:0]; // @[Shift.scala 64:52]
  assign _T_1502 = {_T_1501,1'h0}; // @[Cat.scala 29:58]
  assign _T_1503 = _T_1499 ? _T_1502 : _T_1498; // @[Shift.scala 64:27]
  assign normalFracTmp = _T_1468 ? _T_1503 : 50'h0; // @[Shift.scala 16:10]
  assign _T_1505 = $signed(greaterScale) + $signed(10'sh2); // @[PositFMA.scala 130:36]
  assign _T_1506 = $signed(_T_1505); // @[PositFMA.scala 130:36]
  assign _T_1507 = {1'h1,_T_1463,_T_1466}; // @[Cat.scala 29:58]
  assign _T_1508 = $signed(_T_1507); // @[PositFMA.scala 130:61]
  assign _GEN_20 = {{3{_T_1508[6]}},_T_1508}; // @[PositFMA.scala 130:42]
  assign _T_1510 = $signed(_T_1506) + $signed(_GEN_20); // @[PositFMA.scala 130:42]
  assign sumScale = $signed(_T_1510); // @[PositFMA.scala 130:42]
  assign sumFrac = normalFracTmp[49:26]; // @[PositFMA.scala 131:41]
  assign grsTmp = normalFracTmp[25:0]; // @[PositFMA.scala 134:41]
  assign _T_1511 = grsTmp[25:24]; // @[PositFMA.scala 137:40]
  assign _T_1512 = grsTmp[23:0]; // @[PositFMA.scala 137:56]
  assign _T_1513 = _T_1512 != 24'h0; // @[PositFMA.scala 137:60]
  assign underflow = $signed(sumScale) < $signed(-10'she1); // @[PositFMA.scala 144:32]
  assign overflow = $signed(sumScale) > $signed(10'she0); // @[PositFMA.scala 145:32]
  assign _T_1514 = signSumSig != 52'h0; // @[PositFMA.scala 154:32]
  assign decF_isZero = ~ _T_1514; // @[PositFMA.scala 154:20]
  assign _T_1516 = underflow ? $signed(-10'she1) : $signed(sumScale); // @[Mux.scala 87:16]
  assign _T_1517 = overflow ? $signed(10'she0) : $signed(_T_1516); // @[Mux.scala 87:16]
  assign _GEN_21 = _T_1517[8:0]; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  assign decF_scale = $signed(_GEN_21); // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  assign _T_1518 = decF_scale[2:0]; // @[convert.scala 46:61]
  assign _T_1519 = ~ _T_1518; // @[convert.scala 46:52]
  assign _T_1521 = sumSign ? _T_1519 : _T_1518; // @[convert.scala 46:42]
  assign _T_1522 = decF_scale[8:3]; // @[convert.scala 48:34]
  assign _T_1523 = _T_1522[5:5]; // @[convert.scala 49:36]
  assign _T_1525 = ~ _T_1522; // @[convert.scala 50:36]
  assign _T_1526 = $signed(_T_1525); // @[convert.scala 50:36]
  assign _T_1527 = _T_1523 ? $signed(_T_1526) : $signed(_T_1522); // @[convert.scala 50:28]
  assign _T_1528 = _T_1523 ^ sumSign; // @[convert.scala 51:31]
  assign _T_1529 = ~ _T_1528; // @[convert.scala 52:43]
  assign _T_1533 = {_T_1529,_T_1528,_T_1521,sumFrac,_T_1511,_T_1513}; // @[Cat.scala 29:58]
  assign _T_1534 = $unsigned(_T_1527); // @[Shift.scala 39:17]
  assign _T_1535 = _T_1534 < 6'h20; // @[Shift.scala 39:24]
  assign _T_1536 = _T_1527[4:0]; // @[Shift.scala 40:44]
  assign _T_1537 = _T_1533[31:16]; // @[Shift.scala 90:30]
  assign _T_1538 = _T_1533[15:0]; // @[Shift.scala 90:48]
  assign _T_1539 = _T_1538 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_22 = {{15'd0}, _T_1539}; // @[Shift.scala 90:39]
  assign _T_1540 = _T_1537 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_1541 = _T_1536[4]; // @[Shift.scala 12:21]
  assign _T_1542 = _T_1533[31]; // @[Shift.scala 12:21]
  assign _T_1544 = _T_1542 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_1545 = {_T_1544,_T_1540}; // @[Cat.scala 29:58]
  assign _T_1546 = _T_1541 ? _T_1545 : _T_1533; // @[Shift.scala 91:22]
  assign _T_1547 = _T_1536[3:0]; // @[Shift.scala 92:77]
  assign _T_1548 = _T_1546[31:8]; // @[Shift.scala 90:30]
  assign _T_1549 = _T_1546[7:0]; // @[Shift.scala 90:48]
  assign _T_1550 = _T_1549 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_23 = {{23'd0}, _T_1550}; // @[Shift.scala 90:39]
  assign _T_1551 = _T_1548 | _GEN_23; // @[Shift.scala 90:39]
  assign _T_1552 = _T_1547[3]; // @[Shift.scala 12:21]
  assign _T_1553 = _T_1546[31]; // @[Shift.scala 12:21]
  assign _T_1555 = _T_1553 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_1556 = {_T_1555,_T_1551}; // @[Cat.scala 29:58]
  assign _T_1557 = _T_1552 ? _T_1556 : _T_1546; // @[Shift.scala 91:22]
  assign _T_1558 = _T_1547[2:0]; // @[Shift.scala 92:77]
  assign _T_1559 = _T_1557[31:4]; // @[Shift.scala 90:30]
  assign _T_1560 = _T_1557[3:0]; // @[Shift.scala 90:48]
  assign _T_1561 = _T_1560 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_24 = {{27'd0}, _T_1561}; // @[Shift.scala 90:39]
  assign _T_1562 = _T_1559 | _GEN_24; // @[Shift.scala 90:39]
  assign _T_1563 = _T_1558[2]; // @[Shift.scala 12:21]
  assign _T_1564 = _T_1557[31]; // @[Shift.scala 12:21]
  assign _T_1566 = _T_1564 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_1567 = {_T_1566,_T_1562}; // @[Cat.scala 29:58]
  assign _T_1568 = _T_1563 ? _T_1567 : _T_1557; // @[Shift.scala 91:22]
  assign _T_1569 = _T_1558[1:0]; // @[Shift.scala 92:77]
  assign _T_1570 = _T_1568[31:2]; // @[Shift.scala 90:30]
  assign _T_1571 = _T_1568[1:0]; // @[Shift.scala 90:48]
  assign _T_1572 = _T_1571 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_25 = {{29'd0}, _T_1572}; // @[Shift.scala 90:39]
  assign _T_1573 = _T_1570 | _GEN_25; // @[Shift.scala 90:39]
  assign _T_1574 = _T_1569[1]; // @[Shift.scala 12:21]
  assign _T_1575 = _T_1568[31]; // @[Shift.scala 12:21]
  assign _T_1577 = _T_1575 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_1578 = {_T_1577,_T_1573}; // @[Cat.scala 29:58]
  assign _T_1579 = _T_1574 ? _T_1578 : _T_1568; // @[Shift.scala 91:22]
  assign _T_1580 = _T_1569[0:0]; // @[Shift.scala 92:77]
  assign _T_1581 = _T_1579[31:1]; // @[Shift.scala 90:30]
  assign _T_1582 = _T_1579[0:0]; // @[Shift.scala 90:48]
  assign _GEN_26 = {{30'd0}, _T_1582}; // @[Shift.scala 90:39]
  assign _T_1584 = _T_1581 | _GEN_26; // @[Shift.scala 90:39]
  assign _T_1586 = _T_1579[31]; // @[Shift.scala 12:21]
  assign _T_1587 = {_T_1586,_T_1584}; // @[Cat.scala 29:58]
  assign _T_1588 = _T_1580 ? _T_1587 : _T_1579; // @[Shift.scala 91:22]
  assign _T_1591 = _T_1542 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 71:12]
  assign _T_1592 = _T_1535 ? _T_1588 : _T_1591; // @[Shift.scala 39:10]
  assign _T_1593 = _T_1592[3]; // @[convert.scala 55:31]
  assign _T_1594 = _T_1592[2]; // @[convert.scala 56:31]
  assign _T_1595 = _T_1592[1]; // @[convert.scala 57:31]
  assign _T_1596 = _T_1592[0]; // @[convert.scala 58:31]
  assign _T_1597 = _T_1592[31:3]; // @[convert.scala 59:69]
  assign _T_1598 = _T_1597 != 29'h0; // @[convert.scala 59:81]
  assign _T_1599 = ~ _T_1598; // @[convert.scala 59:50]
  assign _T_1601 = _T_1597 == 29'h1fffffff; // @[convert.scala 60:81]
  assign _T_1602 = _T_1593 | _T_1595; // @[convert.scala 61:44]
  assign _T_1603 = _T_1602 | _T_1596; // @[convert.scala 61:52]
  assign _T_1604 = _T_1594 & _T_1603; // @[convert.scala 61:36]
  assign _T_1605 = ~ _T_1601; // @[convert.scala 62:63]
  assign _T_1606 = _T_1605 & _T_1604; // @[convert.scala 62:103]
  assign _T_1607 = _T_1599 | _T_1606; // @[convert.scala 62:60]
  assign _GEN_27 = {{28'd0}, _T_1607}; // @[convert.scala 63:56]
  assign _T_1610 = _T_1597 + _GEN_27; // @[convert.scala 63:56]
  assign _T_1611 = {sumSign,_T_1610}; // @[Cat.scala 29:58]
  assign io_F = _T_1619; // @[PositFMA.scala 174:15]
  assign io_outValid = _T_1615; // @[PositFMA.scala 173:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  outIsNaR_phase2 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  mulSig_phase2 = _RAND_1[50:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  addFrac_phase2 = _RAND_2[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mulScale_phase2 = _RAND_3[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addScale_phase2 = _RAND_4[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addSign_phase2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addZero_phase2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  inValid_phase2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1615 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_1619 = _RAND_9[29:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (io_inValid) begin
      outIsNaR_phase2 <= outIsNaR;
    end
    if (io_inValid) begin
      mulSig_phase2 <= mulSig;
    end
    if (io_inValid) begin
      addFrac_phase2 <= decC_fraction;
    end
    if (io_inValid) begin
      mulScale_phase2 <= mulScale;
    end
    if (io_inValid) begin
      addScale_phase2 <= decC_scale;
    end
    if (io_inValid) begin
      addSign_phase2 <= _T_601;
    end
    if (io_inValid) begin
      addZero_phase2 <= decC_isZero;
    end
    if (reset) begin
      inValid_phase2 <= 1'h0;
    end else begin
      inValid_phase2 <= io_inValid;
    end
    if (reset) begin
      _T_1615 <= 1'h0;
    end else begin
      _T_1615 <= inValid_phase2;
    end
    if (inValid_phase2) begin
      if (outIsNaR_phase2) begin
        _T_1619 <= 30'h20000000;
      end else begin
        if (decF_isZero) begin
          _T_1619 <= 30'h0;
        end else begin
          _T_1619 <= _T_1611;
        end
      end
    end
  end
endmodule
