module PositDivSqrter16_1(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input  [15:0] io_A,
  input  [15:0] io_B,
  output        io_diviValid,
  output        io_sqrtValid,
  output        io_invalidExc,
  output [15:0] io_Q
);
  reg [4:0] cycleNum; // @[PositDivisionSqrt.scala 63:26]
  reg [31:0] _RAND_0;
  reg  sqrtOp_Z; // @[PositDivisionSqrt.scala 65:22]
  reg [31:0] _RAND_1;
  reg  isNaR_Z; // @[PositDivisionSqrt.scala 66:22]
  reg [31:0] _RAND_2;
  reg  isZero_Z; // @[PositDivisionSqrt.scala 67:22]
  reg [31:0] _RAND_3;
  reg [6:0] scale_Z; // @[PositDivisionSqrt.scala 68:22]
  reg [31:0] _RAND_4;
  reg  signB_Z; // @[PositDivisionSqrt.scala 69:28]
  reg [31:0] _RAND_5;
  reg [11:0] fractB_Z; // @[PositDivisionSqrt.scala 70:22]
  reg [31:0] _RAND_6;
  reg [18:0] rem_Z; // @[PositDivisionSqrt.scala 71:22]
  reg [31:0] _RAND_7;
  reg [18:0] sigX_Z; // @[PositDivisionSqrt.scala 72:22]
  reg [31:0] _RAND_8;
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [13:0] _T_4; // @[convert.scala 19:24]
  wire [13:0] _T_5; // @[convert.scala 19:43]
  wire [13:0] _T_6; // @[convert.scala 19:39]
  wire [7:0] _T_7; // @[LZD.scala 43:32]
  wire [3:0] _T_8; // @[LZD.scala 43:32]
  wire [1:0] _T_9; // @[LZD.scala 43:32]
  wire  _T_10; // @[LZD.scala 39:14]
  wire  _T_11; // @[LZD.scala 39:21]
  wire  _T_12; // @[LZD.scala 39:30]
  wire  _T_13; // @[LZD.scala 39:27]
  wire  _T_14; // @[LZD.scala 39:25]
  wire [1:0] _T_15; // @[Cat.scala 29:58]
  wire [1:0] _T_16; // @[LZD.scala 44:32]
  wire  _T_17; // @[LZD.scala 39:14]
  wire  _T_18; // @[LZD.scala 39:21]
  wire  _T_19; // @[LZD.scala 39:30]
  wire  _T_20; // @[LZD.scala 39:27]
  wire  _T_21; // @[LZD.scala 39:25]
  wire [1:0] _T_22; // @[Cat.scala 29:58]
  wire  _T_23; // @[Shift.scala 12:21]
  wire  _T_24; // @[Shift.scala 12:21]
  wire  _T_25; // @[LZD.scala 49:16]
  wire  _T_26; // @[LZD.scala 49:27]
  wire  _T_27; // @[LZD.scala 49:25]
  wire  _T_28; // @[LZD.scala 49:47]
  wire  _T_29; // @[LZD.scala 49:59]
  wire  _T_30; // @[LZD.scala 49:35]
  wire [2:0] _T_32; // @[Cat.scala 29:58]
  wire [3:0] _T_33; // @[LZD.scala 44:32]
  wire [1:0] _T_34; // @[LZD.scala 43:32]
  wire  _T_35; // @[LZD.scala 39:14]
  wire  _T_36; // @[LZD.scala 39:21]
  wire  _T_37; // @[LZD.scala 39:30]
  wire  _T_38; // @[LZD.scala 39:27]
  wire  _T_39; // @[LZD.scala 39:25]
  wire [1:0] _T_40; // @[Cat.scala 29:58]
  wire [1:0] _T_41; // @[LZD.scala 44:32]
  wire  _T_42; // @[LZD.scala 39:14]
  wire  _T_43; // @[LZD.scala 39:21]
  wire  _T_44; // @[LZD.scala 39:30]
  wire  _T_45; // @[LZD.scala 39:27]
  wire  _T_46; // @[LZD.scala 39:25]
  wire [1:0] _T_47; // @[Cat.scala 29:58]
  wire  _T_48; // @[Shift.scala 12:21]
  wire  _T_49; // @[Shift.scala 12:21]
  wire  _T_50; // @[LZD.scala 49:16]
  wire  _T_51; // @[LZD.scala 49:27]
  wire  _T_52; // @[LZD.scala 49:25]
  wire  _T_53; // @[LZD.scala 49:47]
  wire  _T_54; // @[LZD.scala 49:59]
  wire  _T_55; // @[LZD.scala 49:35]
  wire [2:0] _T_57; // @[Cat.scala 29:58]
  wire  _T_58; // @[Shift.scala 12:21]
  wire  _T_59; // @[Shift.scala 12:21]
  wire  _T_60; // @[LZD.scala 49:16]
  wire  _T_61; // @[LZD.scala 49:27]
  wire  _T_62; // @[LZD.scala 49:25]
  wire [1:0] _T_63; // @[LZD.scala 49:47]
  wire [1:0] _T_64; // @[LZD.scala 49:59]
  wire [1:0] _T_65; // @[LZD.scala 49:35]
  wire [3:0] _T_67; // @[Cat.scala 29:58]
  wire [5:0] _T_68; // @[LZD.scala 44:32]
  wire [3:0] _T_69; // @[LZD.scala 43:32]
  wire [1:0] _T_70; // @[LZD.scala 43:32]
  wire  _T_71; // @[LZD.scala 39:14]
  wire  _T_72; // @[LZD.scala 39:21]
  wire  _T_73; // @[LZD.scala 39:30]
  wire  _T_74; // @[LZD.scala 39:27]
  wire  _T_75; // @[LZD.scala 39:25]
  wire [1:0] _T_76; // @[Cat.scala 29:58]
  wire [1:0] _T_77; // @[LZD.scala 44:32]
  wire  _T_78; // @[LZD.scala 39:14]
  wire  _T_79; // @[LZD.scala 39:21]
  wire  _T_80; // @[LZD.scala 39:30]
  wire  _T_81; // @[LZD.scala 39:27]
  wire  _T_82; // @[LZD.scala 39:25]
  wire [1:0] _T_83; // @[Cat.scala 29:58]
  wire  _T_84; // @[Shift.scala 12:21]
  wire  _T_85; // @[Shift.scala 12:21]
  wire  _T_86; // @[LZD.scala 49:16]
  wire  _T_87; // @[LZD.scala 49:27]
  wire  _T_88; // @[LZD.scala 49:25]
  wire  _T_89; // @[LZD.scala 49:47]
  wire  _T_90; // @[LZD.scala 49:59]
  wire  _T_91; // @[LZD.scala 49:35]
  wire [2:0] _T_93; // @[Cat.scala 29:58]
  wire [1:0] _T_94; // @[LZD.scala 44:32]
  wire  _T_95; // @[LZD.scala 39:14]
  wire  _T_96; // @[LZD.scala 39:21]
  wire  _T_97; // @[LZD.scala 39:30]
  wire  _T_98; // @[LZD.scala 39:27]
  wire  _T_99; // @[LZD.scala 39:25]
  wire [1:0] _T_100; // @[Cat.scala 29:58]
  wire  _T_101; // @[Shift.scala 12:21]
  wire [1:0] _T_103; // @[LZD.scala 55:32]
  wire [1:0] _T_104; // @[LZD.scala 55:20]
  wire [2:0] _T_105; // @[Cat.scala 29:58]
  wire  _T_106; // @[Shift.scala 12:21]
  wire [2:0] _T_108; // @[LZD.scala 55:32]
  wire [2:0] _T_109; // @[LZD.scala 55:20]
  wire [3:0] _T_110; // @[Cat.scala 29:58]
  wire [3:0] _T_111; // @[convert.scala 21:22]
  wire [12:0] _T_112; // @[convert.scala 22:36]
  wire  _T_113; // @[Shift.scala 16:24]
  wire  _T_115; // @[Shift.scala 12:21]
  wire [4:0] _T_116; // @[Shift.scala 64:52]
  wire [12:0] _T_118; // @[Cat.scala 29:58]
  wire [12:0] _T_119; // @[Shift.scala 64:27]
  wire [2:0] _T_120; // @[Shift.scala 66:70]
  wire  _T_121; // @[Shift.scala 12:21]
  wire [8:0] _T_122; // @[Shift.scala 64:52]
  wire [12:0] _T_124; // @[Cat.scala 29:58]
  wire [12:0] _T_125; // @[Shift.scala 64:27]
  wire [1:0] _T_126; // @[Shift.scala 66:70]
  wire  _T_127; // @[Shift.scala 12:21]
  wire [10:0] _T_128; // @[Shift.scala 64:52]
  wire [12:0] _T_130; // @[Cat.scala 29:58]
  wire [12:0] _T_131; // @[Shift.scala 64:27]
  wire  _T_132; // @[Shift.scala 66:70]
  wire [11:0] _T_134; // @[Shift.scala 64:52]
  wire [12:0] _T_135; // @[Cat.scala 29:58]
  wire [12:0] _T_136; // @[Shift.scala 64:27]
  wire [12:0] _T_137; // @[Shift.scala 16:10]
  wire  _T_138; // @[convert.scala 23:34]
  wire [11:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_140; // @[convert.scala 25:26]
  wire [3:0] _T_142; // @[convert.scala 25:42]
  wire  _T_145; // @[convert.scala 26:67]
  wire  _T_146; // @[convert.scala 26:51]
  wire [5:0] _T_147; // @[Cat.scala 29:58]
  wire [14:0] _T_149; // @[convert.scala 29:56]
  wire  _T_150; // @[convert.scala 29:60]
  wire  _T_151; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_154; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [5:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_163; // @[convert.scala 18:24]
  wire  _T_164; // @[convert.scala 18:40]
  wire  _T_165; // @[convert.scala 18:36]
  wire [13:0] _T_166; // @[convert.scala 19:24]
  wire [13:0] _T_167; // @[convert.scala 19:43]
  wire [13:0] _T_168; // @[convert.scala 19:39]
  wire [7:0] _T_169; // @[LZD.scala 43:32]
  wire [3:0] _T_170; // @[LZD.scala 43:32]
  wire [1:0] _T_171; // @[LZD.scala 43:32]
  wire  _T_172; // @[LZD.scala 39:14]
  wire  _T_173; // @[LZD.scala 39:21]
  wire  _T_174; // @[LZD.scala 39:30]
  wire  _T_175; // @[LZD.scala 39:27]
  wire  _T_176; // @[LZD.scala 39:25]
  wire [1:0] _T_177; // @[Cat.scala 29:58]
  wire [1:0] _T_178; // @[LZD.scala 44:32]
  wire  _T_179; // @[LZD.scala 39:14]
  wire  _T_180; // @[LZD.scala 39:21]
  wire  _T_181; // @[LZD.scala 39:30]
  wire  _T_182; // @[LZD.scala 39:27]
  wire  _T_183; // @[LZD.scala 39:25]
  wire [1:0] _T_184; // @[Cat.scala 29:58]
  wire  _T_185; // @[Shift.scala 12:21]
  wire  _T_186; // @[Shift.scala 12:21]
  wire  _T_187; // @[LZD.scala 49:16]
  wire  _T_188; // @[LZD.scala 49:27]
  wire  _T_189; // @[LZD.scala 49:25]
  wire  _T_190; // @[LZD.scala 49:47]
  wire  _T_191; // @[LZD.scala 49:59]
  wire  _T_192; // @[LZD.scala 49:35]
  wire [2:0] _T_194; // @[Cat.scala 29:58]
  wire [3:0] _T_195; // @[LZD.scala 44:32]
  wire [1:0] _T_196; // @[LZD.scala 43:32]
  wire  _T_197; // @[LZD.scala 39:14]
  wire  _T_198; // @[LZD.scala 39:21]
  wire  _T_199; // @[LZD.scala 39:30]
  wire  _T_200; // @[LZD.scala 39:27]
  wire  _T_201; // @[LZD.scala 39:25]
  wire [1:0] _T_202; // @[Cat.scala 29:58]
  wire [1:0] _T_203; // @[LZD.scala 44:32]
  wire  _T_204; // @[LZD.scala 39:14]
  wire  _T_205; // @[LZD.scala 39:21]
  wire  _T_206; // @[LZD.scala 39:30]
  wire  _T_207; // @[LZD.scala 39:27]
  wire  _T_208; // @[LZD.scala 39:25]
  wire [1:0] _T_209; // @[Cat.scala 29:58]
  wire  _T_210; // @[Shift.scala 12:21]
  wire  _T_211; // @[Shift.scala 12:21]
  wire  _T_212; // @[LZD.scala 49:16]
  wire  _T_213; // @[LZD.scala 49:27]
  wire  _T_214; // @[LZD.scala 49:25]
  wire  _T_215; // @[LZD.scala 49:47]
  wire  _T_216; // @[LZD.scala 49:59]
  wire  _T_217; // @[LZD.scala 49:35]
  wire [2:0] _T_219; // @[Cat.scala 29:58]
  wire  _T_220; // @[Shift.scala 12:21]
  wire  _T_221; // @[Shift.scala 12:21]
  wire  _T_222; // @[LZD.scala 49:16]
  wire  _T_223; // @[LZD.scala 49:27]
  wire  _T_224; // @[LZD.scala 49:25]
  wire [1:0] _T_225; // @[LZD.scala 49:47]
  wire [1:0] _T_226; // @[LZD.scala 49:59]
  wire [1:0] _T_227; // @[LZD.scala 49:35]
  wire [3:0] _T_229; // @[Cat.scala 29:58]
  wire [5:0] _T_230; // @[LZD.scala 44:32]
  wire [3:0] _T_231; // @[LZD.scala 43:32]
  wire [1:0] _T_232; // @[LZD.scala 43:32]
  wire  _T_233; // @[LZD.scala 39:14]
  wire  _T_234; // @[LZD.scala 39:21]
  wire  _T_235; // @[LZD.scala 39:30]
  wire  _T_236; // @[LZD.scala 39:27]
  wire  _T_237; // @[LZD.scala 39:25]
  wire [1:0] _T_238; // @[Cat.scala 29:58]
  wire [1:0] _T_239; // @[LZD.scala 44:32]
  wire  _T_240; // @[LZD.scala 39:14]
  wire  _T_241; // @[LZD.scala 39:21]
  wire  _T_242; // @[LZD.scala 39:30]
  wire  _T_243; // @[LZD.scala 39:27]
  wire  _T_244; // @[LZD.scala 39:25]
  wire [1:0] _T_245; // @[Cat.scala 29:58]
  wire  _T_246; // @[Shift.scala 12:21]
  wire  _T_247; // @[Shift.scala 12:21]
  wire  _T_248; // @[LZD.scala 49:16]
  wire  _T_249; // @[LZD.scala 49:27]
  wire  _T_250; // @[LZD.scala 49:25]
  wire  _T_251; // @[LZD.scala 49:47]
  wire  _T_252; // @[LZD.scala 49:59]
  wire  _T_253; // @[LZD.scala 49:35]
  wire [2:0] _T_255; // @[Cat.scala 29:58]
  wire [1:0] _T_256; // @[LZD.scala 44:32]
  wire  _T_257; // @[LZD.scala 39:14]
  wire  _T_258; // @[LZD.scala 39:21]
  wire  _T_259; // @[LZD.scala 39:30]
  wire  _T_260; // @[LZD.scala 39:27]
  wire  _T_261; // @[LZD.scala 39:25]
  wire [1:0] _T_262; // @[Cat.scala 29:58]
  wire  _T_263; // @[Shift.scala 12:21]
  wire [1:0] _T_265; // @[LZD.scala 55:32]
  wire [1:0] _T_266; // @[LZD.scala 55:20]
  wire [2:0] _T_267; // @[Cat.scala 29:58]
  wire  _T_268; // @[Shift.scala 12:21]
  wire [2:0] _T_270; // @[LZD.scala 55:32]
  wire [2:0] _T_271; // @[LZD.scala 55:20]
  wire [3:0] _T_272; // @[Cat.scala 29:58]
  wire [3:0] _T_273; // @[convert.scala 21:22]
  wire [12:0] _T_274; // @[convert.scala 22:36]
  wire  _T_275; // @[Shift.scala 16:24]
  wire  _T_277; // @[Shift.scala 12:21]
  wire [4:0] _T_278; // @[Shift.scala 64:52]
  wire [12:0] _T_280; // @[Cat.scala 29:58]
  wire [12:0] _T_281; // @[Shift.scala 64:27]
  wire [2:0] _T_282; // @[Shift.scala 66:70]
  wire  _T_283; // @[Shift.scala 12:21]
  wire [8:0] _T_284; // @[Shift.scala 64:52]
  wire [12:0] _T_286; // @[Cat.scala 29:58]
  wire [12:0] _T_287; // @[Shift.scala 64:27]
  wire [1:0] _T_288; // @[Shift.scala 66:70]
  wire  _T_289; // @[Shift.scala 12:21]
  wire [10:0] _T_290; // @[Shift.scala 64:52]
  wire [12:0] _T_292; // @[Cat.scala 29:58]
  wire [12:0] _T_293; // @[Shift.scala 64:27]
  wire  _T_294; // @[Shift.scala 66:70]
  wire [11:0] _T_296; // @[Shift.scala 64:52]
  wire [12:0] _T_297; // @[Cat.scala 29:58]
  wire [12:0] _T_298; // @[Shift.scala 64:27]
  wire [12:0] _T_299; // @[Shift.scala 16:10]
  wire  _T_300; // @[convert.scala 23:34]
  wire [11:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_302; // @[convert.scala 25:26]
  wire [3:0] _T_304; // @[convert.scala 25:42]
  wire  _T_307; // @[convert.scala 26:67]
  wire  _T_308; // @[convert.scala 26:51]
  wire [5:0] _T_309; // @[Cat.scala 29:58]
  wire [14:0] _T_311; // @[convert.scala 29:56]
  wire  _T_312; // @[convert.scala 29:60]
  wire  _T_313; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_316; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [5:0] decB_scale; // @[convert.scala 32:24]
  wire [2:0] _T_325; // @[Bitwise.scala 71:12]
  wire  _T_326; // @[PositDivisionSqrt.scala 80:40]
  wire [18:0] sigA_S; // @[Cat.scala 29:58]
  wire  _T_329; // @[PositDivisionSqrt.scala 82:31]
  wire [18:0] sigB_S; // @[Cat.scala 29:58]
  wire  _T_332; // @[PositDivisionSqrt.scala 85:25]
  wire  invalidSqrt; // @[PositDivisionSqrt.scala 85:37]
  wire  _T_333; // @[PositDivisionSqrt.scala 88:42]
  wire  _T_334; // @[PositDivisionSqrt.scala 89:42]
  wire  _T_335; // @[PositDivisionSqrt.scala 89:56]
  wire  _T_336; // @[PositDivisionSqrt.scala 94:46]
  wire  _T_337; // @[PositDivisionSqrt.scala 94:43]
  wire  _T_338; // @[PositDivisionSqrt.scala 94:62]
  wire  _T_339; // @[PositDivisionSqrt.scala 94:59]
  wire  specialCaseA_S; // @[PositDivisionSqrt.scala 97:38]
  wire  specialCaseB_S; // @[PositDivisionSqrt.scala 98:38]
  wire  _T_340; // @[PositDivisionSqrt.scala 99:27]
  wire  _T_341; // @[PositDivisionSqrt.scala 99:46]
  wire  normalCase_S_div; // @[PositDivisionSqrt.scala 99:43]
  wire  normalCase_S_sqrt; // @[PositDivisionSqrt.scala 100:43]
  wire  normalCase_S; // @[PositDivisionSqrt.scala 101:30]
  wire [6:0] sExpQuot_S_div; // @[PositDivisionSqrt.scala 103:38]
  wire  _T_344; // @[PositDivisionSqrt.scala 104:50]
  wire  oddSqrt_S; // @[PositDivisionSqrt.scala 104:37]
  wire  idle; // @[PositDivisionSqrt.scala 109:39]
  wire  ready; // @[PositDivisionSqrt.scala 110:39]
  wire  entering; // @[PositDivisionSqrt.scala 111:35]
  wire  entering_normalCase; // @[PositDivisionSqrt.scala 112:38]
  wire  _T_345; // @[PositDivisionSqrt.scala 113:35]
  wire  _T_346; // @[PositDivisionSqrt.scala 113:58]
  wire  scaleNotChange; // @[PositDivisionSqrt.scala 113:50]
  wire  _T_347; // @[PositDivisionSqrt.scala 114:39]
  wire  skipCycle2; // @[PositDivisionSqrt.scala 114:48]
  wire  _T_348; // @[PositDivisionSqrt.scala 116:8]
  wire  _T_349; // @[PositDivisionSqrt.scala 116:14]
  wire  _T_350; // @[PositDivisionSqrt.scala 117:32]
  wire  _T_351; // @[PositDivisionSqrt.scala 117:30]
  wire [4:0] _T_353; // @[PositDivisionSqrt.scala 119:26]
  wire [4:0] _T_354; // @[PositDivisionSqrt.scala 118:20]
  wire [4:0] _GEN_9; // @[PositDivisionSqrt.scala 117:64]
  wire [4:0] _T_355; // @[PositDivisionSqrt.scala 117:64]
  wire  _T_357; // @[PositDivisionSqrt.scala 123:30]
  wire  _T_358; // @[PositDivisionSqrt.scala 123:27]
  wire [4:0] _T_360; // @[PositDivisionSqrt.scala 123:52]
  wire [4:0] _T_361; // @[PositDivisionSqrt.scala 123:20]
  wire [4:0] _T_362; // @[PositDivisionSqrt.scala 122:64]
  wire  _T_364; // @[PositDivisionSqrt.scala 124:27]
  wire [4:0] _GEN_10; // @[PositDivisionSqrt.scala 123:64]
  wire [4:0] _T_366; // @[PositDivisionSqrt.scala 123:64]
  wire [4:0] _T_367; // @[PositDivisionSqrt.scala 134:42]
  wire  _T_369; // @[PositDivisionSqrt.scala 137:31]
  wire  _T_370; // @[PositDivisionSqrt.scala 137:28]
  wire [31:0] _T_371; // @[PositDivisionSqrt.scala 146:22]
  wire [29:0] _T_372; // @[PositDivisionSqrt.scala 146:35]
  wire  _T_373; // @[PositDivisionSqrt.scala 148:26]
  wire  _T_374; // @[PositDivisionSqrt.scala 148:23]
  wire [18:0] _T_375; // @[PositDivisionSqrt.scala 148:16]
  wire  _T_376; // @[PositDivisionSqrt.scala 149:23]
  wire [19:0] _T_377; // @[PositDivisionSqrt.scala 149:46]
  wire [18:0] _T_378; // @[PositDivisionSqrt.scala 149:56]
  wire [18:0] _T_379; // @[PositDivisionSqrt.scala 149:16]
  wire [18:0] _T_380; // @[PositDivisionSqrt.scala 148:66]
  wire  _T_381; // @[PositDivisionSqrt.scala 150:17]
  wire [18:0] _T_382; // @[PositDivisionSqrt.scala 150:16]
  wire [18:0] rem; // @[PositDivisionSqrt.scala 149:66]
  wire  _T_384; // @[PositDivisionSqrt.scala 152:29]
  wire [18:0] _T_385; // @[PositDivisionSqrt.scala 152:22]
  wire  _T_386; // @[PositDivisionSqrt.scala 153:29]
  wire [15:0] _T_387; // @[PositDivisionSqrt.scala 153:22]
  wire [18:0] _GEN_11; // @[PositDivisionSqrt.scala 152:93]
  wire [18:0] _T_388; // @[PositDivisionSqrt.scala 152:93]
  wire  _T_390; // @[PositDivisionSqrt.scala 154:33]
  wire  _T_391; // @[PositDivisionSqrt.scala 154:30]
  wire  _T_392; // @[PositDivisionSqrt.scala 154:57]
  wire [18:0] _T_395; // @[Cat.scala 29:58]
  wire [18:0] _T_396; // @[PositDivisionSqrt.scala 154:22]
  wire [18:0] _T_397; // @[PositDivisionSqrt.scala 153:93]
  wire  _T_399; // @[PositDivisionSqrt.scala 155:30]
  wire  _T_400; // @[PositDivisionSqrt.scala 156:83]
  wire [14:0] _T_402; // @[Bitwise.scala 71:12]
  wire [17:0] bitMask; // @[PositDivisionSqrt.scala 145:21 PositDivisionSqrt.scala 146:14]
  wire [17:0] _GEN_12; // @[PositDivisionSqrt.scala 156:53]
  wire [17:0] _T_403; // @[PositDivisionSqrt.scala 156:53]
  wire [18:0] _GEN_13; // @[PositDivisionSqrt.scala 155:51]
  wire [18:0] _T_404; // @[PositDivisionSqrt.scala 155:51]
  wire [16:0] _T_405; // @[PositDivisionSqrt.scala 157:53]
  wire [18:0] _GEN_14; // @[PositDivisionSqrt.scala 156:89]
  wire [18:0] _T_406; // @[PositDivisionSqrt.scala 156:89]
  wire [18:0] _T_407; // @[PositDivisionSqrt.scala 155:22]
  wire [18:0] trialTerm; // @[PositDivisionSqrt.scala 154:93]
  wire  _T_409; // @[PositDivisionSqrt.scala 162:56]
  wire  _T_410; // @[PositDivisionSqrt.scala 162:40]
  wire [18:0] _T_413; // @[PositDivisionSqrt.scala 163:97]
  wire [18:0] _T_415; // @[PositDivisionSqrt.scala 164:97]
  wire [18:0] _T_416; // @[PositDivisionSqrt.scala 161:92]
  wire [19:0] _T_421; // @[PositDivisionSqrt.scala 168:98]
  wire [18:0] _T_422; // @[PositDivisionSqrt.scala 168:108]
  wire [18:0] _T_424; // @[PositDivisionSqrt.scala 168:112]
  wire [18:0] _T_428; // @[PositDivisionSqrt.scala 169:112]
  wire [18:0] _T_429; // @[PositDivisionSqrt.scala 166:26]
  wire [18:0] trialRem; // @[PositDivisionSqrt.scala 159:27]
  wire  _T_430; // @[PositDivisionSqrt.scala 173:35]
  wire  trIsZero; // @[PositDivisionSqrt.scala 173:25]
  wire  _T_431; // @[PositDivisionSqrt.scala 174:30]
  wire  remIsZero; // @[PositDivisionSqrt.scala 174:25]
  wire  _T_433; // @[PositDivisionSqrt.scala 176:64]
  wire  _T_434; // @[PositDivisionSqrt.scala 176:49]
  wire  _T_435; // @[PositDivisionSqrt.scala 176:29]
  wire  _T_436; // @[PositDivisionSqrt.scala 178:61]
  wire  _T_437; // @[PositDivisionSqrt.scala 178:49]
  wire  _T_439; // @[Mux.scala 87:16]
  wire  newBit; // @[Mux.scala 87:16]
  wire  _T_440; // @[PositDivisionSqrt.scala 183:41]
  wire  _T_441; // @[PositDivisionSqrt.scala 183:51]
  wire  _T_442; // @[PositDivisionSqrt.scala 183:48]
  wire  _T_443; // @[PositDivisionSqrt.scala 183:28]
  wire  _T_446; // @[PositDivisionSqrt.scala 187:39]
  wire  _T_447; // @[PositDivisionSqrt.scala 187:28]
  wire [18:0] _T_450; // @[PositDivisionSqrt.scala 188:47]
  wire [18:0] _T_451; // @[PositDivisionSqrt.scala 188:18]
  wire [16:0] _T_453; // @[PositDivisionSqrt.scala 189:18]
  wire [18:0] _GEN_15; // @[PositDivisionSqrt.scala 188:78]
  wire [18:0] _T_454; // @[PositDivisionSqrt.scala 188:78]
  wire [18:0] _GEN_16; // @[PositDivisionSqrt.scala 190:47]
  wire [18:0] _T_456; // @[PositDivisionSqrt.scala 190:47]
  wire [18:0] _T_457; // @[PositDivisionSqrt.scala 190:18]
  wire [18:0] _T_458; // @[PositDivisionSqrt.scala 189:78]
  wire [1:0] _T_460; // @[PositDivisionSqrt.scala 196:53]
  wire [1:0] sigXBias; // @[PositDivisionSqrt.scala 196:21]
  wire [18:0] _GEN_17; // @[PositDivisionSqrt.scala 197:25]
  wire [18:0] realSigX; // @[PositDivisionSqrt.scala 197:25]
  wire [11:0] _T_463; // @[PositDivisionSqrt.scala 200:97]
  wire [11:0] _T_464; // @[PositDivisionSqrt.scala 201:97]
  wire [11:0] realFrac; // @[PositDivisionSqrt.scala 198:21]
  wire  _T_465; // @[PositDivisionSqrt.scala 205:33]
  wire  _T_466; // @[PositDivisionSqrt.scala 205:58]
  wire  _T_467; // @[PositDivisionSqrt.scala 205:48]
  wire  scaleNeedSub; // @[PositDivisionSqrt.scala 205:23]
  wire  _T_469; // @[PositDivisionSqrt.scala 206:56]
  wire  notNeedSubTwo; // @[PositDivisionSqrt.scala 206:46]
  wire  scaleSubOne; // @[PositDivisionSqrt.scala 207:36]
  wire  _T_470; // @[PositDivisionSqrt.scala 208:38]
  wire  scaleSubTwo; // @[PositDivisionSqrt.scala 208:36]
  wire [1:0] _T_471; // @[Cat.scala 29:58]
  wire [2:0] _T_472; // @[PositDivisionSqrt.scala 209:63]
  wire [6:0] _GEN_18; // @[PositDivisionSqrt.scala 209:31]
  wire [6:0] _T_474; // @[PositDivisionSqrt.scala 209:31]
  wire [6:0] realExp; // @[PositDivisionSqrt.scala 209:31]
  wire  underflow; // @[PositDivisionSqrt.scala 210:31]
  wire  overflow; // @[PositDivisionSqrt.scala 211:31]
  wire  decQ_sign; // @[PositDivisionSqrt.scala 215:33]
  wire [6:0] _T_476; // @[Mux.scala 87:16]
  wire [6:0] _T_477; // @[Mux.scala 87:16]
  wire [2:0] _T_478; // @[PositDivisionSqrt.scala 224:48]
  wire [2:0] _T_479; // @[PositDivisionSqrt.scala 224:64]
  wire [2:0] decQ_grs; // @[PositDivisionSqrt.scala 224:23]
  wire  outValid; // @[PositDivisionSqrt.scala 229:28]
  wire [5:0] _GEN_19; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire [5:0] decQ_scale; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire  _T_485; // @[convert.scala 46:61]
  wire  _T_486; // @[convert.scala 46:52]
  wire  _T_488; // @[convert.scala 46:42]
  wire [4:0] _T_489; // @[convert.scala 48:34]
  wire  _T_490; // @[convert.scala 49:36]
  wire [4:0] _T_492; // @[convert.scala 50:36]
  wire [4:0] _T_493; // @[convert.scala 50:36]
  wire [4:0] _T_494; // @[convert.scala 50:28]
  wire  _T_495; // @[convert.scala 51:31]
  wire  _T_496; // @[convert.scala 52:43]
  wire [17:0] _T_500; // @[Cat.scala 29:58]
  wire [4:0] _T_501; // @[Shift.scala 39:17]
  wire  _T_502; // @[Shift.scala 39:24]
  wire [1:0] _T_504; // @[Shift.scala 90:30]
  wire [15:0] _T_505; // @[Shift.scala 90:48]
  wire  _T_506; // @[Shift.scala 90:57]
  wire [1:0] _GEN_20; // @[Shift.scala 90:39]
  wire [1:0] _T_507; // @[Shift.scala 90:39]
  wire  _T_508; // @[Shift.scala 12:21]
  wire  _T_509; // @[Shift.scala 12:21]
  wire [15:0] _T_511; // @[Bitwise.scala 71:12]
  wire [17:0] _T_512; // @[Cat.scala 29:58]
  wire [17:0] _T_513; // @[Shift.scala 91:22]
  wire [3:0] _T_514; // @[Shift.scala 92:77]
  wire [9:0] _T_515; // @[Shift.scala 90:30]
  wire [7:0] _T_516; // @[Shift.scala 90:48]
  wire  _T_517; // @[Shift.scala 90:57]
  wire [9:0] _GEN_21; // @[Shift.scala 90:39]
  wire [9:0] _T_518; // @[Shift.scala 90:39]
  wire  _T_519; // @[Shift.scala 12:21]
  wire  _T_520; // @[Shift.scala 12:21]
  wire [7:0] _T_522; // @[Bitwise.scala 71:12]
  wire [17:0] _T_523; // @[Cat.scala 29:58]
  wire [17:0] _T_524; // @[Shift.scala 91:22]
  wire [2:0] _T_525; // @[Shift.scala 92:77]
  wire [13:0] _T_526; // @[Shift.scala 90:30]
  wire [3:0] _T_527; // @[Shift.scala 90:48]
  wire  _T_528; // @[Shift.scala 90:57]
  wire [13:0] _GEN_22; // @[Shift.scala 90:39]
  wire [13:0] _T_529; // @[Shift.scala 90:39]
  wire  _T_530; // @[Shift.scala 12:21]
  wire  _T_531; // @[Shift.scala 12:21]
  wire [3:0] _T_533; // @[Bitwise.scala 71:12]
  wire [17:0] _T_534; // @[Cat.scala 29:58]
  wire [17:0] _T_535; // @[Shift.scala 91:22]
  wire [1:0] _T_536; // @[Shift.scala 92:77]
  wire [15:0] _T_537; // @[Shift.scala 90:30]
  wire [1:0] _T_538; // @[Shift.scala 90:48]
  wire  _T_539; // @[Shift.scala 90:57]
  wire [15:0] _GEN_23; // @[Shift.scala 90:39]
  wire [15:0] _T_540; // @[Shift.scala 90:39]
  wire  _T_541; // @[Shift.scala 12:21]
  wire  _T_542; // @[Shift.scala 12:21]
  wire [1:0] _T_544; // @[Bitwise.scala 71:12]
  wire [17:0] _T_545; // @[Cat.scala 29:58]
  wire [17:0] _T_546; // @[Shift.scala 91:22]
  wire  _T_547; // @[Shift.scala 92:77]
  wire [16:0] _T_548; // @[Shift.scala 90:30]
  wire  _T_549; // @[Shift.scala 90:48]
  wire [16:0] _GEN_24; // @[Shift.scala 90:39]
  wire [16:0] _T_551; // @[Shift.scala 90:39]
  wire  _T_553; // @[Shift.scala 12:21]
  wire [17:0] _T_554; // @[Cat.scala 29:58]
  wire [17:0] _T_555; // @[Shift.scala 91:22]
  wire [17:0] _T_558; // @[Bitwise.scala 71:12]
  wire [17:0] _T_559; // @[Shift.scala 39:10]
  wire  _T_560; // @[convert.scala 55:31]
  wire  _T_561; // @[convert.scala 56:31]
  wire  _T_562; // @[convert.scala 57:31]
  wire  _T_563; // @[convert.scala 58:31]
  wire [14:0] _T_564; // @[convert.scala 59:69]
  wire  _T_565; // @[convert.scala 59:81]
  wire  _T_566; // @[convert.scala 59:50]
  wire  _T_568; // @[convert.scala 60:81]
  wire  _T_569; // @[convert.scala 61:44]
  wire  _T_570; // @[convert.scala 61:52]
  wire  _T_571; // @[convert.scala 61:36]
  wire  _T_572; // @[convert.scala 62:63]
  wire  _T_573; // @[convert.scala 62:103]
  wire  _T_574; // @[convert.scala 62:60]
  wire [14:0] _GEN_25; // @[convert.scala 63:56]
  wire [14:0] _T_577; // @[convert.scala 63:56]
  wire [15:0] _T_578; // @[Cat.scala 29:58]
  wire [15:0] _T_580; // @[Mux.scala 87:16]
  assign _T_1 = io_A[15]; // @[convert.scala 18:24]
  assign _T_2 = io_A[14]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[14:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[13:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[13:6]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[7:4]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8[3:2]; // @[LZD.scala 43:32]
  assign _T_10 = _T_9 != 2'h0; // @[LZD.scala 39:14]
  assign _T_11 = _T_9[1]; // @[LZD.scala 39:21]
  assign _T_12 = _T_9[0]; // @[LZD.scala 39:30]
  assign _T_13 = ~ _T_12; // @[LZD.scala 39:27]
  assign _T_14 = _T_11 | _T_13; // @[LZD.scala 39:25]
  assign _T_15 = {_T_10,_T_14}; // @[Cat.scala 29:58]
  assign _T_16 = _T_8[1:0]; // @[LZD.scala 44:32]
  assign _T_17 = _T_16 != 2'h0; // @[LZD.scala 39:14]
  assign _T_18 = _T_16[1]; // @[LZD.scala 39:21]
  assign _T_19 = _T_16[0]; // @[LZD.scala 39:30]
  assign _T_20 = ~ _T_19; // @[LZD.scala 39:27]
  assign _T_21 = _T_18 | _T_20; // @[LZD.scala 39:25]
  assign _T_22 = {_T_17,_T_21}; // @[Cat.scala 29:58]
  assign _T_23 = _T_15[1]; // @[Shift.scala 12:21]
  assign _T_24 = _T_22[1]; // @[Shift.scala 12:21]
  assign _T_25 = _T_23 | _T_24; // @[LZD.scala 49:16]
  assign _T_26 = ~ _T_24; // @[LZD.scala 49:27]
  assign _T_27 = _T_23 | _T_26; // @[LZD.scala 49:25]
  assign _T_28 = _T_15[0:0]; // @[LZD.scala 49:47]
  assign _T_29 = _T_22[0:0]; // @[LZD.scala 49:59]
  assign _T_30 = _T_23 ? _T_28 : _T_29; // @[LZD.scala 49:35]
  assign _T_32 = {_T_25,_T_27,_T_30}; // @[Cat.scala 29:58]
  assign _T_33 = _T_7[3:0]; // @[LZD.scala 44:32]
  assign _T_34 = _T_33[3:2]; // @[LZD.scala 43:32]
  assign _T_35 = _T_34 != 2'h0; // @[LZD.scala 39:14]
  assign _T_36 = _T_34[1]; // @[LZD.scala 39:21]
  assign _T_37 = _T_34[0]; // @[LZD.scala 39:30]
  assign _T_38 = ~ _T_37; // @[LZD.scala 39:27]
  assign _T_39 = _T_36 | _T_38; // @[LZD.scala 39:25]
  assign _T_40 = {_T_35,_T_39}; // @[Cat.scala 29:58]
  assign _T_41 = _T_33[1:0]; // @[LZD.scala 44:32]
  assign _T_42 = _T_41 != 2'h0; // @[LZD.scala 39:14]
  assign _T_43 = _T_41[1]; // @[LZD.scala 39:21]
  assign _T_44 = _T_41[0]; // @[LZD.scala 39:30]
  assign _T_45 = ~ _T_44; // @[LZD.scala 39:27]
  assign _T_46 = _T_43 | _T_45; // @[LZD.scala 39:25]
  assign _T_47 = {_T_42,_T_46}; // @[Cat.scala 29:58]
  assign _T_48 = _T_40[1]; // @[Shift.scala 12:21]
  assign _T_49 = _T_47[1]; // @[Shift.scala 12:21]
  assign _T_50 = _T_48 | _T_49; // @[LZD.scala 49:16]
  assign _T_51 = ~ _T_49; // @[LZD.scala 49:27]
  assign _T_52 = _T_48 | _T_51; // @[LZD.scala 49:25]
  assign _T_53 = _T_40[0:0]; // @[LZD.scala 49:47]
  assign _T_54 = _T_47[0:0]; // @[LZD.scala 49:59]
  assign _T_55 = _T_48 ? _T_53 : _T_54; // @[LZD.scala 49:35]
  assign _T_57 = {_T_50,_T_52,_T_55}; // @[Cat.scala 29:58]
  assign _T_58 = _T_32[2]; // @[Shift.scala 12:21]
  assign _T_59 = _T_57[2]; // @[Shift.scala 12:21]
  assign _T_60 = _T_58 | _T_59; // @[LZD.scala 49:16]
  assign _T_61 = ~ _T_59; // @[LZD.scala 49:27]
  assign _T_62 = _T_58 | _T_61; // @[LZD.scala 49:25]
  assign _T_63 = _T_32[1:0]; // @[LZD.scala 49:47]
  assign _T_64 = _T_57[1:0]; // @[LZD.scala 49:59]
  assign _T_65 = _T_58 ? _T_63 : _T_64; // @[LZD.scala 49:35]
  assign _T_67 = {_T_60,_T_62,_T_65}; // @[Cat.scala 29:58]
  assign _T_68 = _T_6[5:0]; // @[LZD.scala 44:32]
  assign _T_69 = _T_68[5:2]; // @[LZD.scala 43:32]
  assign _T_70 = _T_69[3:2]; // @[LZD.scala 43:32]
  assign _T_71 = _T_70 != 2'h0; // @[LZD.scala 39:14]
  assign _T_72 = _T_70[1]; // @[LZD.scala 39:21]
  assign _T_73 = _T_70[0]; // @[LZD.scala 39:30]
  assign _T_74 = ~ _T_73; // @[LZD.scala 39:27]
  assign _T_75 = _T_72 | _T_74; // @[LZD.scala 39:25]
  assign _T_76 = {_T_71,_T_75}; // @[Cat.scala 29:58]
  assign _T_77 = _T_69[1:0]; // @[LZD.scala 44:32]
  assign _T_78 = _T_77 != 2'h0; // @[LZD.scala 39:14]
  assign _T_79 = _T_77[1]; // @[LZD.scala 39:21]
  assign _T_80 = _T_77[0]; // @[LZD.scala 39:30]
  assign _T_81 = ~ _T_80; // @[LZD.scala 39:27]
  assign _T_82 = _T_79 | _T_81; // @[LZD.scala 39:25]
  assign _T_83 = {_T_78,_T_82}; // @[Cat.scala 29:58]
  assign _T_84 = _T_76[1]; // @[Shift.scala 12:21]
  assign _T_85 = _T_83[1]; // @[Shift.scala 12:21]
  assign _T_86 = _T_84 | _T_85; // @[LZD.scala 49:16]
  assign _T_87 = ~ _T_85; // @[LZD.scala 49:27]
  assign _T_88 = _T_84 | _T_87; // @[LZD.scala 49:25]
  assign _T_89 = _T_76[0:0]; // @[LZD.scala 49:47]
  assign _T_90 = _T_83[0:0]; // @[LZD.scala 49:59]
  assign _T_91 = _T_84 ? _T_89 : _T_90; // @[LZD.scala 49:35]
  assign _T_93 = {_T_86,_T_88,_T_91}; // @[Cat.scala 29:58]
  assign _T_94 = _T_68[1:0]; // @[LZD.scala 44:32]
  assign _T_95 = _T_94 != 2'h0; // @[LZD.scala 39:14]
  assign _T_96 = _T_94[1]; // @[LZD.scala 39:21]
  assign _T_97 = _T_94[0]; // @[LZD.scala 39:30]
  assign _T_98 = ~ _T_97; // @[LZD.scala 39:27]
  assign _T_99 = _T_96 | _T_98; // @[LZD.scala 39:25]
  assign _T_100 = {_T_95,_T_99}; // @[Cat.scala 29:58]
  assign _T_101 = _T_93[2]; // @[Shift.scala 12:21]
  assign _T_103 = _T_93[1:0]; // @[LZD.scala 55:32]
  assign _T_104 = _T_101 ? _T_103 : _T_100; // @[LZD.scala 55:20]
  assign _T_105 = {_T_101,_T_104}; // @[Cat.scala 29:58]
  assign _T_106 = _T_67[3]; // @[Shift.scala 12:21]
  assign _T_108 = _T_67[2:0]; // @[LZD.scala 55:32]
  assign _T_109 = _T_106 ? _T_108 : _T_105; // @[LZD.scala 55:20]
  assign _T_110 = {_T_106,_T_109}; // @[Cat.scala 29:58]
  assign _T_111 = ~ _T_110; // @[convert.scala 21:22]
  assign _T_112 = io_A[12:0]; // @[convert.scala 22:36]
  assign _T_113 = _T_111 < 4'hd; // @[Shift.scala 16:24]
  assign _T_115 = _T_111[3]; // @[Shift.scala 12:21]
  assign _T_116 = _T_112[4:0]; // @[Shift.scala 64:52]
  assign _T_118 = {_T_116,8'h0}; // @[Cat.scala 29:58]
  assign _T_119 = _T_115 ? _T_118 : _T_112; // @[Shift.scala 64:27]
  assign _T_120 = _T_111[2:0]; // @[Shift.scala 66:70]
  assign _T_121 = _T_120[2]; // @[Shift.scala 12:21]
  assign _T_122 = _T_119[8:0]; // @[Shift.scala 64:52]
  assign _T_124 = {_T_122,4'h0}; // @[Cat.scala 29:58]
  assign _T_125 = _T_121 ? _T_124 : _T_119; // @[Shift.scala 64:27]
  assign _T_126 = _T_120[1:0]; // @[Shift.scala 66:70]
  assign _T_127 = _T_126[1]; // @[Shift.scala 12:21]
  assign _T_128 = _T_125[10:0]; // @[Shift.scala 64:52]
  assign _T_130 = {_T_128,2'h0}; // @[Cat.scala 29:58]
  assign _T_131 = _T_127 ? _T_130 : _T_125; // @[Shift.scala 64:27]
  assign _T_132 = _T_126[0:0]; // @[Shift.scala 66:70]
  assign _T_134 = _T_131[11:0]; // @[Shift.scala 64:52]
  assign _T_135 = {_T_134,1'h0}; // @[Cat.scala 29:58]
  assign _T_136 = _T_132 ? _T_135 : _T_131; // @[Shift.scala 64:27]
  assign _T_137 = _T_113 ? _T_136 : 13'h0; // @[Shift.scala 16:10]
  assign _T_138 = _T_137[12:12]; // @[convert.scala 23:34]
  assign decA_fraction = _T_137[11:0]; // @[convert.scala 24:34]
  assign _T_140 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_142 = _T_3 ? _T_111 : _T_110; // @[convert.scala 25:42]
  assign _T_145 = ~ _T_138; // @[convert.scala 26:67]
  assign _T_146 = _T_1 ? _T_145 : _T_138; // @[convert.scala 26:51]
  assign _T_147 = {_T_140,_T_142,_T_146}; // @[Cat.scala 29:58]
  assign _T_149 = io_A[14:0]; // @[convert.scala 29:56]
  assign _T_150 = _T_149 != 15'h0; // @[convert.scala 29:60]
  assign _T_151 = ~ _T_150; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_151; // @[convert.scala 29:39]
  assign _T_154 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_154 & _T_151; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_147); // @[convert.scala 32:24]
  assign _T_163 = io_B[15]; // @[convert.scala 18:24]
  assign _T_164 = io_B[14]; // @[convert.scala 18:40]
  assign _T_165 = _T_163 ^ _T_164; // @[convert.scala 18:36]
  assign _T_166 = io_B[14:1]; // @[convert.scala 19:24]
  assign _T_167 = io_B[13:0]; // @[convert.scala 19:43]
  assign _T_168 = _T_166 ^ _T_167; // @[convert.scala 19:39]
  assign _T_169 = _T_168[13:6]; // @[LZD.scala 43:32]
  assign _T_170 = _T_169[7:4]; // @[LZD.scala 43:32]
  assign _T_171 = _T_170[3:2]; // @[LZD.scala 43:32]
  assign _T_172 = _T_171 != 2'h0; // @[LZD.scala 39:14]
  assign _T_173 = _T_171[1]; // @[LZD.scala 39:21]
  assign _T_174 = _T_171[0]; // @[LZD.scala 39:30]
  assign _T_175 = ~ _T_174; // @[LZD.scala 39:27]
  assign _T_176 = _T_173 | _T_175; // @[LZD.scala 39:25]
  assign _T_177 = {_T_172,_T_176}; // @[Cat.scala 29:58]
  assign _T_178 = _T_170[1:0]; // @[LZD.scala 44:32]
  assign _T_179 = _T_178 != 2'h0; // @[LZD.scala 39:14]
  assign _T_180 = _T_178[1]; // @[LZD.scala 39:21]
  assign _T_181 = _T_178[0]; // @[LZD.scala 39:30]
  assign _T_182 = ~ _T_181; // @[LZD.scala 39:27]
  assign _T_183 = _T_180 | _T_182; // @[LZD.scala 39:25]
  assign _T_184 = {_T_179,_T_183}; // @[Cat.scala 29:58]
  assign _T_185 = _T_177[1]; // @[Shift.scala 12:21]
  assign _T_186 = _T_184[1]; // @[Shift.scala 12:21]
  assign _T_187 = _T_185 | _T_186; // @[LZD.scala 49:16]
  assign _T_188 = ~ _T_186; // @[LZD.scala 49:27]
  assign _T_189 = _T_185 | _T_188; // @[LZD.scala 49:25]
  assign _T_190 = _T_177[0:0]; // @[LZD.scala 49:47]
  assign _T_191 = _T_184[0:0]; // @[LZD.scala 49:59]
  assign _T_192 = _T_185 ? _T_190 : _T_191; // @[LZD.scala 49:35]
  assign _T_194 = {_T_187,_T_189,_T_192}; // @[Cat.scala 29:58]
  assign _T_195 = _T_169[3:0]; // @[LZD.scala 44:32]
  assign _T_196 = _T_195[3:2]; // @[LZD.scala 43:32]
  assign _T_197 = _T_196 != 2'h0; // @[LZD.scala 39:14]
  assign _T_198 = _T_196[1]; // @[LZD.scala 39:21]
  assign _T_199 = _T_196[0]; // @[LZD.scala 39:30]
  assign _T_200 = ~ _T_199; // @[LZD.scala 39:27]
  assign _T_201 = _T_198 | _T_200; // @[LZD.scala 39:25]
  assign _T_202 = {_T_197,_T_201}; // @[Cat.scala 29:58]
  assign _T_203 = _T_195[1:0]; // @[LZD.scala 44:32]
  assign _T_204 = _T_203 != 2'h0; // @[LZD.scala 39:14]
  assign _T_205 = _T_203[1]; // @[LZD.scala 39:21]
  assign _T_206 = _T_203[0]; // @[LZD.scala 39:30]
  assign _T_207 = ~ _T_206; // @[LZD.scala 39:27]
  assign _T_208 = _T_205 | _T_207; // @[LZD.scala 39:25]
  assign _T_209 = {_T_204,_T_208}; // @[Cat.scala 29:58]
  assign _T_210 = _T_202[1]; // @[Shift.scala 12:21]
  assign _T_211 = _T_209[1]; // @[Shift.scala 12:21]
  assign _T_212 = _T_210 | _T_211; // @[LZD.scala 49:16]
  assign _T_213 = ~ _T_211; // @[LZD.scala 49:27]
  assign _T_214 = _T_210 | _T_213; // @[LZD.scala 49:25]
  assign _T_215 = _T_202[0:0]; // @[LZD.scala 49:47]
  assign _T_216 = _T_209[0:0]; // @[LZD.scala 49:59]
  assign _T_217 = _T_210 ? _T_215 : _T_216; // @[LZD.scala 49:35]
  assign _T_219 = {_T_212,_T_214,_T_217}; // @[Cat.scala 29:58]
  assign _T_220 = _T_194[2]; // @[Shift.scala 12:21]
  assign _T_221 = _T_219[2]; // @[Shift.scala 12:21]
  assign _T_222 = _T_220 | _T_221; // @[LZD.scala 49:16]
  assign _T_223 = ~ _T_221; // @[LZD.scala 49:27]
  assign _T_224 = _T_220 | _T_223; // @[LZD.scala 49:25]
  assign _T_225 = _T_194[1:0]; // @[LZD.scala 49:47]
  assign _T_226 = _T_219[1:0]; // @[LZD.scala 49:59]
  assign _T_227 = _T_220 ? _T_225 : _T_226; // @[LZD.scala 49:35]
  assign _T_229 = {_T_222,_T_224,_T_227}; // @[Cat.scala 29:58]
  assign _T_230 = _T_168[5:0]; // @[LZD.scala 44:32]
  assign _T_231 = _T_230[5:2]; // @[LZD.scala 43:32]
  assign _T_232 = _T_231[3:2]; // @[LZD.scala 43:32]
  assign _T_233 = _T_232 != 2'h0; // @[LZD.scala 39:14]
  assign _T_234 = _T_232[1]; // @[LZD.scala 39:21]
  assign _T_235 = _T_232[0]; // @[LZD.scala 39:30]
  assign _T_236 = ~ _T_235; // @[LZD.scala 39:27]
  assign _T_237 = _T_234 | _T_236; // @[LZD.scala 39:25]
  assign _T_238 = {_T_233,_T_237}; // @[Cat.scala 29:58]
  assign _T_239 = _T_231[1:0]; // @[LZD.scala 44:32]
  assign _T_240 = _T_239 != 2'h0; // @[LZD.scala 39:14]
  assign _T_241 = _T_239[1]; // @[LZD.scala 39:21]
  assign _T_242 = _T_239[0]; // @[LZD.scala 39:30]
  assign _T_243 = ~ _T_242; // @[LZD.scala 39:27]
  assign _T_244 = _T_241 | _T_243; // @[LZD.scala 39:25]
  assign _T_245 = {_T_240,_T_244}; // @[Cat.scala 29:58]
  assign _T_246 = _T_238[1]; // @[Shift.scala 12:21]
  assign _T_247 = _T_245[1]; // @[Shift.scala 12:21]
  assign _T_248 = _T_246 | _T_247; // @[LZD.scala 49:16]
  assign _T_249 = ~ _T_247; // @[LZD.scala 49:27]
  assign _T_250 = _T_246 | _T_249; // @[LZD.scala 49:25]
  assign _T_251 = _T_238[0:0]; // @[LZD.scala 49:47]
  assign _T_252 = _T_245[0:0]; // @[LZD.scala 49:59]
  assign _T_253 = _T_246 ? _T_251 : _T_252; // @[LZD.scala 49:35]
  assign _T_255 = {_T_248,_T_250,_T_253}; // @[Cat.scala 29:58]
  assign _T_256 = _T_230[1:0]; // @[LZD.scala 44:32]
  assign _T_257 = _T_256 != 2'h0; // @[LZD.scala 39:14]
  assign _T_258 = _T_256[1]; // @[LZD.scala 39:21]
  assign _T_259 = _T_256[0]; // @[LZD.scala 39:30]
  assign _T_260 = ~ _T_259; // @[LZD.scala 39:27]
  assign _T_261 = _T_258 | _T_260; // @[LZD.scala 39:25]
  assign _T_262 = {_T_257,_T_261}; // @[Cat.scala 29:58]
  assign _T_263 = _T_255[2]; // @[Shift.scala 12:21]
  assign _T_265 = _T_255[1:0]; // @[LZD.scala 55:32]
  assign _T_266 = _T_263 ? _T_265 : _T_262; // @[LZD.scala 55:20]
  assign _T_267 = {_T_263,_T_266}; // @[Cat.scala 29:58]
  assign _T_268 = _T_229[3]; // @[Shift.scala 12:21]
  assign _T_270 = _T_229[2:0]; // @[LZD.scala 55:32]
  assign _T_271 = _T_268 ? _T_270 : _T_267; // @[LZD.scala 55:20]
  assign _T_272 = {_T_268,_T_271}; // @[Cat.scala 29:58]
  assign _T_273 = ~ _T_272; // @[convert.scala 21:22]
  assign _T_274 = io_B[12:0]; // @[convert.scala 22:36]
  assign _T_275 = _T_273 < 4'hd; // @[Shift.scala 16:24]
  assign _T_277 = _T_273[3]; // @[Shift.scala 12:21]
  assign _T_278 = _T_274[4:0]; // @[Shift.scala 64:52]
  assign _T_280 = {_T_278,8'h0}; // @[Cat.scala 29:58]
  assign _T_281 = _T_277 ? _T_280 : _T_274; // @[Shift.scala 64:27]
  assign _T_282 = _T_273[2:0]; // @[Shift.scala 66:70]
  assign _T_283 = _T_282[2]; // @[Shift.scala 12:21]
  assign _T_284 = _T_281[8:0]; // @[Shift.scala 64:52]
  assign _T_286 = {_T_284,4'h0}; // @[Cat.scala 29:58]
  assign _T_287 = _T_283 ? _T_286 : _T_281; // @[Shift.scala 64:27]
  assign _T_288 = _T_282[1:0]; // @[Shift.scala 66:70]
  assign _T_289 = _T_288[1]; // @[Shift.scala 12:21]
  assign _T_290 = _T_287[10:0]; // @[Shift.scala 64:52]
  assign _T_292 = {_T_290,2'h0}; // @[Cat.scala 29:58]
  assign _T_293 = _T_289 ? _T_292 : _T_287; // @[Shift.scala 64:27]
  assign _T_294 = _T_288[0:0]; // @[Shift.scala 66:70]
  assign _T_296 = _T_293[11:0]; // @[Shift.scala 64:52]
  assign _T_297 = {_T_296,1'h0}; // @[Cat.scala 29:58]
  assign _T_298 = _T_294 ? _T_297 : _T_293; // @[Shift.scala 64:27]
  assign _T_299 = _T_275 ? _T_298 : 13'h0; // @[Shift.scala 16:10]
  assign _T_300 = _T_299[12:12]; // @[convert.scala 23:34]
  assign decB_fraction = _T_299[11:0]; // @[convert.scala 24:34]
  assign _T_302 = _T_165 == 1'h0; // @[convert.scala 25:26]
  assign _T_304 = _T_165 ? _T_273 : _T_272; // @[convert.scala 25:42]
  assign _T_307 = ~ _T_300; // @[convert.scala 26:67]
  assign _T_308 = _T_163 ? _T_307 : _T_300; // @[convert.scala 26:51]
  assign _T_309 = {_T_302,_T_304,_T_308}; // @[Cat.scala 29:58]
  assign _T_311 = io_B[14:0]; // @[convert.scala 29:56]
  assign _T_312 = _T_311 != 15'h0; // @[convert.scala 29:60]
  assign _T_313 = ~ _T_312; // @[convert.scala 29:41]
  assign decB_isNaR = _T_163 & _T_313; // @[convert.scala 29:39]
  assign _T_316 = _T_163 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_316 & _T_313; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_309); // @[convert.scala 32:24]
  assign _T_325 = _T_1 ? 3'h7 : 3'h0; // @[Bitwise.scala 71:12]
  assign _T_326 = ~ _T_1; // @[PositDivisionSqrt.scala 80:40]
  assign sigA_S = {_T_325,_T_326,decA_fraction,3'h0}; // @[Cat.scala 29:58]
  assign _T_329 = ~ _T_163; // @[PositDivisionSqrt.scala 82:31]
  assign sigB_S = {_T_163,_T_329,decB_fraction,5'h0}; // @[Cat.scala 29:58]
  assign _T_332 = decA_isNaR == 1'h0; // @[PositDivisionSqrt.scala 85:25]
  assign invalidSqrt = _T_332 & _T_1; // @[PositDivisionSqrt.scala 85:37]
  assign _T_333 = decA_isNaR | invalidSqrt; // @[PositDivisionSqrt.scala 88:42]
  assign _T_334 = decA_isNaR | decB_isNaR; // @[PositDivisionSqrt.scala 89:42]
  assign _T_335 = _T_334 | decB_isZero; // @[PositDivisionSqrt.scala 89:56]
  assign _T_336 = decB_isZero == 1'h0; // @[PositDivisionSqrt.scala 94:46]
  assign _T_337 = decA_isZero & _T_336; // @[PositDivisionSqrt.scala 94:43]
  assign _T_338 = decB_isNaR == 1'h0; // @[PositDivisionSqrt.scala 94:62]
  assign _T_339 = _T_337 & _T_338; // @[PositDivisionSqrt.scala 94:59]
  assign specialCaseA_S = decA_isNaR | decA_isZero; // @[PositDivisionSqrt.scala 97:38]
  assign specialCaseB_S = decB_isNaR | decB_isZero; // @[PositDivisionSqrt.scala 98:38]
  assign _T_340 = specialCaseA_S == 1'h0; // @[PositDivisionSqrt.scala 99:27]
  assign _T_341 = specialCaseB_S == 1'h0; // @[PositDivisionSqrt.scala 99:46]
  assign normalCase_S_div = _T_340 & _T_341; // @[PositDivisionSqrt.scala 99:43]
  assign normalCase_S_sqrt = _T_340 & _T_154; // @[PositDivisionSqrt.scala 100:43]
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div; // @[PositDivisionSqrt.scala 101:30]
  assign sExpQuot_S_div = $signed(decA_scale) - $signed(decB_scale); // @[PositDivisionSqrt.scala 103:38]
  assign _T_344 = decA_scale[0]; // @[PositDivisionSqrt.scala 104:50]
  assign oddSqrt_S = io_sqrtOp & _T_344; // @[PositDivisionSqrt.scala 104:37]
  assign idle = cycleNum == 5'h0; // @[PositDivisionSqrt.scala 109:39]
  assign ready = cycleNum <= 5'h1; // @[PositDivisionSqrt.scala 110:39]
  assign entering = ready & io_inValid; // @[PositDivisionSqrt.scala 111:35]
  assign entering_normalCase = entering & normalCase_S; // @[PositDivisionSqrt.scala 112:38]
  assign _T_345 = sigX_Z[18]; // @[PositDivisionSqrt.scala 113:35]
  assign _T_346 = sigX_Z[16]; // @[PositDivisionSqrt.scala 113:58]
  assign scaleNotChange = _T_345 ^ _T_346; // @[PositDivisionSqrt.scala 113:50]
  assign _T_347 = cycleNum == 5'h3; // @[PositDivisionSqrt.scala 114:39]
  assign skipCycle2 = _T_347 & scaleNotChange; // @[PositDivisionSqrt.scala 114:48]
  assign _T_348 = idle == 1'h0; // @[PositDivisionSqrt.scala 116:8]
  assign _T_349 = _T_348 | io_inValid; // @[PositDivisionSqrt.scala 116:14]
  assign _T_350 = normalCase_S == 1'h0; // @[PositDivisionSqrt.scala 117:32]
  assign _T_351 = entering & _T_350; // @[PositDivisionSqrt.scala 117:30]
  assign _T_353 = io_sqrtOp ? 5'h11 : 5'h13; // @[PositDivisionSqrt.scala 119:26]
  assign _T_354 = entering_normalCase ? _T_353 : 5'h0; // @[PositDivisionSqrt.scala 118:20]
  assign _GEN_9 = {{4'd0}, _T_351}; // @[PositDivisionSqrt.scala 117:64]
  assign _T_355 = _GEN_9 | _T_354; // @[PositDivisionSqrt.scala 117:64]
  assign _T_357 = skipCycle2 == 1'h0; // @[PositDivisionSqrt.scala 123:30]
  assign _T_358 = _T_348 & _T_357; // @[PositDivisionSqrt.scala 123:27]
  assign _T_360 = cycleNum - 5'h1; // @[PositDivisionSqrt.scala 123:52]
  assign _T_361 = _T_358 ? _T_360 : 5'h0; // @[PositDivisionSqrt.scala 123:20]
  assign _T_362 = _T_355 | _T_361; // @[PositDivisionSqrt.scala 122:64]
  assign _T_364 = _T_348 & skipCycle2; // @[PositDivisionSqrt.scala 124:27]
  assign _GEN_10 = {{4'd0}, _T_364}; // @[PositDivisionSqrt.scala 123:64]
  assign _T_366 = _T_362 | _GEN_10; // @[PositDivisionSqrt.scala 123:64]
  assign _T_367 = decA_scale[5:1]; // @[PositDivisionSqrt.scala 134:42]
  assign _T_369 = io_sqrtOp == 1'h0; // @[PositDivisionSqrt.scala 137:31]
  assign _T_370 = entering_normalCase & _T_369; // @[PositDivisionSqrt.scala 137:28]
  assign _T_371 = 32'h1 << cycleNum; // @[PositDivisionSqrt.scala 146:22]
  assign _T_372 = _T_371[31:2]; // @[PositDivisionSqrt.scala 146:35]
  assign _T_373 = oddSqrt_S == 1'h0; // @[PositDivisionSqrt.scala 148:26]
  assign _T_374 = ready & _T_373; // @[PositDivisionSqrt.scala 148:23]
  assign _T_375 = _T_374 ? sigA_S : 19'h0; // @[PositDivisionSqrt.scala 148:16]
  assign _T_376 = ready & oddSqrt_S; // @[PositDivisionSqrt.scala 149:23]
  assign _T_377 = {sigA_S, 1'h0}; // @[PositDivisionSqrt.scala 149:46]
  assign _T_378 = _T_377[18:0]; // @[PositDivisionSqrt.scala 149:56]
  assign _T_379 = _T_376 ? _T_378 : 19'h0; // @[PositDivisionSqrt.scala 149:16]
  assign _T_380 = _T_375 | _T_379; // @[PositDivisionSqrt.scala 148:66]
  assign _T_381 = ready == 1'h0; // @[PositDivisionSqrt.scala 150:17]
  assign _T_382 = _T_381 ? rem_Z : 19'h0; // @[PositDivisionSqrt.scala 150:16]
  assign rem = _T_380 | _T_382; // @[PositDivisionSqrt.scala 149:66]
  assign _T_384 = ready & _T_369; // @[PositDivisionSqrt.scala 152:29]
  assign _T_385 = _T_384 ? sigB_S : 19'h0; // @[PositDivisionSqrt.scala 152:22]
  assign _T_386 = ready & io_sqrtOp; // @[PositDivisionSqrt.scala 153:29]
  assign _T_387 = _T_386 ? 16'h8000 : 16'h0; // @[PositDivisionSqrt.scala 153:22]
  assign _GEN_11 = {{3'd0}, _T_387}; // @[PositDivisionSqrt.scala 152:93]
  assign _T_388 = _T_385 | _GEN_11; // @[PositDivisionSqrt.scala 152:93]
  assign _T_390 = sqrtOp_Z == 1'h0; // @[PositDivisionSqrt.scala 154:33]
  assign _T_391 = _T_381 & _T_390; // @[PositDivisionSqrt.scala 154:30]
  assign _T_392 = ~ signB_Z; // @[PositDivisionSqrt.scala 154:57]
  assign _T_395 = {signB_Z,_T_392,fractB_Z,5'h0}; // @[Cat.scala 29:58]
  assign _T_396 = _T_391 ? _T_395 : 19'h0; // @[PositDivisionSqrt.scala 154:22]
  assign _T_397 = _T_388 | _T_396; // @[PositDivisionSqrt.scala 153:93]
  assign _T_399 = _T_381 & sqrtOp_Z; // @[PositDivisionSqrt.scala 155:30]
  assign _T_400 = rem[18:18]; // @[PositDivisionSqrt.scala 156:83]
  assign _T_402 = _T_400 ? 15'h7fff : 15'h0; // @[Bitwise.scala 71:12]
  assign bitMask = _T_372[17:0]; // @[PositDivisionSqrt.scala 145:21 PositDivisionSqrt.scala 146:14]
  assign _GEN_12 = {{3'd0}, _T_402}; // @[PositDivisionSqrt.scala 156:53]
  assign _T_403 = bitMask & _GEN_12; // @[PositDivisionSqrt.scala 156:53]
  assign _GEN_13 = {{1'd0}, _T_403}; // @[PositDivisionSqrt.scala 155:51]
  assign _T_404 = sigX_Z | _GEN_13; // @[PositDivisionSqrt.scala 155:51]
  assign _T_405 = bitMask[17:1]; // @[PositDivisionSqrt.scala 157:53]
  assign _GEN_14 = {{2'd0}, _T_405}; // @[PositDivisionSqrt.scala 156:89]
  assign _T_406 = _T_404 | _GEN_14; // @[PositDivisionSqrt.scala 156:89]
  assign _T_407 = _T_399 ? _T_406 : 19'h0; // @[PositDivisionSqrt.scala 155:22]
  assign trialTerm = _T_397 | _T_407; // @[PositDivisionSqrt.scala 154:93]
  assign _T_409 = trialTerm[18:18]; // @[PositDivisionSqrt.scala 162:56]
  assign _T_410 = _T_400 ^ _T_409; // @[PositDivisionSqrt.scala 162:40]
  assign _T_413 = rem + trialTerm; // @[PositDivisionSqrt.scala 163:97]
  assign _T_415 = rem - trialTerm; // @[PositDivisionSqrt.scala 164:97]
  assign _T_416 = _T_410 ? _T_413 : _T_415; // @[PositDivisionSqrt.scala 161:92]
  assign _T_421 = {rem, 1'h0}; // @[PositDivisionSqrt.scala 168:98]
  assign _T_422 = _T_421[18:0]; // @[PositDivisionSqrt.scala 168:108]
  assign _T_424 = _T_422 + trialTerm; // @[PositDivisionSqrt.scala 168:112]
  assign _T_428 = _T_422 - trialTerm; // @[PositDivisionSqrt.scala 169:112]
  assign _T_429 = _T_410 ? _T_424 : _T_428; // @[PositDivisionSqrt.scala 166:26]
  assign trialRem = ready ? _T_416 : _T_429; // @[PositDivisionSqrt.scala 159:27]
  assign _T_430 = trialRem != 19'h0; // @[PositDivisionSqrt.scala 173:35]
  assign trIsZero = _T_430 == 1'h0; // @[PositDivisionSqrt.scala 173:25]
  assign _T_431 = rem != 19'h0; // @[PositDivisionSqrt.scala 174:30]
  assign remIsZero = _T_431 == 1'h0; // @[PositDivisionSqrt.scala 174:25]
  assign _T_433 = trialRem[18:18]; // @[PositDivisionSqrt.scala 176:64]
  assign _T_434 = _T_409 ^ _T_433; // @[PositDivisionSqrt.scala 176:49]
  assign _T_435 = ~ _T_434; // @[PositDivisionSqrt.scala 176:29]
  assign _T_436 = sigX_Z[18:18]; // @[PositDivisionSqrt.scala 178:61]
  assign _T_437 = ~ _T_436; // @[PositDivisionSqrt.scala 178:49]
  assign _T_439 = remIsZero ? _T_436 : _T_435; // @[Mux.scala 87:16]
  assign newBit = trIsZero ? _T_437 : _T_439; // @[Mux.scala 87:16]
  assign _T_440 = cycleNum > 5'h2; // @[PositDivisionSqrt.scala 183:41]
  assign _T_441 = remIsZero == 1'h0; // @[PositDivisionSqrt.scala 183:51]
  assign _T_442 = _T_440 & _T_441; // @[PositDivisionSqrt.scala 183:48]
  assign _T_443 = entering_normalCase | _T_442; // @[PositDivisionSqrt.scala 183:28]
  assign _T_446 = _T_381 & newBit; // @[PositDivisionSqrt.scala 187:39]
  assign _T_447 = entering_normalCase | _T_446; // @[PositDivisionSqrt.scala 187:28]
  assign _T_450 = {newBit, 18'h0}; // @[PositDivisionSqrt.scala 188:47]
  assign _T_451 = _T_384 ? _T_450 : 19'h0; // @[PositDivisionSqrt.scala 188:18]
  assign _T_453 = _T_386 ? 17'h10000 : 17'h0; // @[PositDivisionSqrt.scala 189:18]
  assign _GEN_15 = {{2'd0}, _T_453}; // @[PositDivisionSqrt.scala 188:78]
  assign _T_454 = _T_451 | _GEN_15; // @[PositDivisionSqrt.scala 188:78]
  assign _GEN_16 = {{1'd0}, bitMask}; // @[PositDivisionSqrt.scala 190:47]
  assign _T_456 = sigX_Z | _GEN_16; // @[PositDivisionSqrt.scala 190:47]
  assign _T_457 = _T_381 ? _T_456 : 19'h0; // @[PositDivisionSqrt.scala 190:18]
  assign _T_458 = _T_454 | _T_457; // @[PositDivisionSqrt.scala 189:78]
  assign _T_460 = {_T_436, 1'h0}; // @[PositDivisionSqrt.scala 196:53]
  assign sigXBias = scaleNotChange ? _T_460 : {{1'd0}, _T_436}; // @[PositDivisionSqrt.scala 196:21]
  assign _GEN_17 = {{17'd0}, sigXBias}; // @[PositDivisionSqrt.scala 197:25]
  assign realSigX = sigX_Z + _GEN_17; // @[PositDivisionSqrt.scala 197:25]
  assign _T_463 = realSigX[15:4]; // @[PositDivisionSqrt.scala 200:97]
  assign _T_464 = realSigX[14:3]; // @[PositDivisionSqrt.scala 201:97]
  assign realFrac = scaleNotChange ? _T_463 : _T_464; // @[PositDivisionSqrt.scala 198:21]
  assign _T_465 = realSigX[18]; // @[PositDivisionSqrt.scala 205:33]
  assign _T_466 = realSigX[16]; // @[PositDivisionSqrt.scala 205:58]
  assign _T_467 = _T_465 ^ _T_466; // @[PositDivisionSqrt.scala 205:48]
  assign scaleNeedSub = ~ _T_467; // @[PositDivisionSqrt.scala 205:23]
  assign _T_469 = realSigX[15]; // @[PositDivisionSqrt.scala 206:56]
  assign notNeedSubTwo = _T_465 ^ _T_469; // @[PositDivisionSqrt.scala 206:46]
  assign scaleSubOne = scaleNeedSub & notNeedSubTwo; // @[PositDivisionSqrt.scala 207:36]
  assign _T_470 = ~ notNeedSubTwo; // @[PositDivisionSqrt.scala 208:38]
  assign scaleSubTwo = scaleNeedSub & _T_470; // @[PositDivisionSqrt.scala 208:36]
  assign _T_471 = {scaleSubTwo,scaleSubOne}; // @[Cat.scala 29:58]
  assign _T_472 = {1'b0,$signed(_T_471)}; // @[PositDivisionSqrt.scala 209:63]
  assign _GEN_18 = {{4{_T_472[2]}},_T_472}; // @[PositDivisionSqrt.scala 209:31]
  assign _T_474 = $signed(scale_Z) - $signed(_GEN_18); // @[PositDivisionSqrt.scala 209:31]
  assign realExp = $signed(_T_474); // @[PositDivisionSqrt.scala 209:31]
  assign underflow = $signed(realExp) < $signed(-7'sh1d); // @[PositDivisionSqrt.scala 210:31]
  assign overflow = $signed(realExp) > $signed(7'sh1c); // @[PositDivisionSqrt.scala 211:31]
  assign decQ_sign = realSigX[18:18]; // @[PositDivisionSqrt.scala 215:33]
  assign _T_476 = underflow ? $signed(-7'sh1d) : $signed(realExp); // @[Mux.scala 87:16]
  assign _T_477 = overflow ? $signed(7'sh1c) : $signed(_T_476); // @[Mux.scala 87:16]
  assign _T_478 = realSigX[3:1]; // @[PositDivisionSqrt.scala 224:48]
  assign _T_479 = realSigX[2:0]; // @[PositDivisionSqrt.scala 224:64]
  assign decQ_grs = scaleNotChange ? _T_478 : _T_479; // @[PositDivisionSqrt.scala 224:23]
  assign outValid = cycleNum == 5'h1; // @[PositDivisionSqrt.scala 229:28]
  assign _GEN_19 = _T_477[5:0]; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign decQ_scale = $signed(_GEN_19); // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign _T_485 = decQ_scale[0]; // @[convert.scala 46:61]
  assign _T_486 = ~ _T_485; // @[convert.scala 46:52]
  assign _T_488 = decQ_sign ? _T_486 : _T_485; // @[convert.scala 46:42]
  assign _T_489 = decQ_scale[5:1]; // @[convert.scala 48:34]
  assign _T_490 = _T_489[4:4]; // @[convert.scala 49:36]
  assign _T_492 = ~ _T_489; // @[convert.scala 50:36]
  assign _T_493 = $signed(_T_492); // @[convert.scala 50:36]
  assign _T_494 = _T_490 ? $signed(_T_493) : $signed(_T_489); // @[convert.scala 50:28]
  assign _T_495 = _T_490 ^ decQ_sign; // @[convert.scala 51:31]
  assign _T_496 = ~ _T_495; // @[convert.scala 52:43]
  assign _T_500 = {_T_496,_T_495,_T_488,realFrac,decQ_grs}; // @[Cat.scala 29:58]
  assign _T_501 = $unsigned(_T_494); // @[Shift.scala 39:17]
  assign _T_502 = _T_501 < 5'h12; // @[Shift.scala 39:24]
  assign _T_504 = _T_500[17:16]; // @[Shift.scala 90:30]
  assign _T_505 = _T_500[15:0]; // @[Shift.scala 90:48]
  assign _T_506 = _T_505 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_20 = {{1'd0}, _T_506}; // @[Shift.scala 90:39]
  assign _T_507 = _T_504 | _GEN_20; // @[Shift.scala 90:39]
  assign _T_508 = _T_501[4]; // @[Shift.scala 12:21]
  assign _T_509 = _T_500[17]; // @[Shift.scala 12:21]
  assign _T_511 = _T_509 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_512 = {_T_511,_T_507}; // @[Cat.scala 29:58]
  assign _T_513 = _T_508 ? _T_512 : _T_500; // @[Shift.scala 91:22]
  assign _T_514 = _T_501[3:0]; // @[Shift.scala 92:77]
  assign _T_515 = _T_513[17:8]; // @[Shift.scala 90:30]
  assign _T_516 = _T_513[7:0]; // @[Shift.scala 90:48]
  assign _T_517 = _T_516 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_21 = {{9'd0}, _T_517}; // @[Shift.scala 90:39]
  assign _T_518 = _T_515 | _GEN_21; // @[Shift.scala 90:39]
  assign _T_519 = _T_514[3]; // @[Shift.scala 12:21]
  assign _T_520 = _T_513[17]; // @[Shift.scala 12:21]
  assign _T_522 = _T_520 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_523 = {_T_522,_T_518}; // @[Cat.scala 29:58]
  assign _T_524 = _T_519 ? _T_523 : _T_513; // @[Shift.scala 91:22]
  assign _T_525 = _T_514[2:0]; // @[Shift.scala 92:77]
  assign _T_526 = _T_524[17:4]; // @[Shift.scala 90:30]
  assign _T_527 = _T_524[3:0]; // @[Shift.scala 90:48]
  assign _T_528 = _T_527 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_22 = {{13'd0}, _T_528}; // @[Shift.scala 90:39]
  assign _T_529 = _T_526 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_530 = _T_525[2]; // @[Shift.scala 12:21]
  assign _T_531 = _T_524[17]; // @[Shift.scala 12:21]
  assign _T_533 = _T_531 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_534 = {_T_533,_T_529}; // @[Cat.scala 29:58]
  assign _T_535 = _T_530 ? _T_534 : _T_524; // @[Shift.scala 91:22]
  assign _T_536 = _T_525[1:0]; // @[Shift.scala 92:77]
  assign _T_537 = _T_535[17:2]; // @[Shift.scala 90:30]
  assign _T_538 = _T_535[1:0]; // @[Shift.scala 90:48]
  assign _T_539 = _T_538 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_23 = {{15'd0}, _T_539}; // @[Shift.scala 90:39]
  assign _T_540 = _T_537 | _GEN_23; // @[Shift.scala 90:39]
  assign _T_541 = _T_536[1]; // @[Shift.scala 12:21]
  assign _T_542 = _T_535[17]; // @[Shift.scala 12:21]
  assign _T_544 = _T_542 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_545 = {_T_544,_T_540}; // @[Cat.scala 29:58]
  assign _T_546 = _T_541 ? _T_545 : _T_535; // @[Shift.scala 91:22]
  assign _T_547 = _T_536[0:0]; // @[Shift.scala 92:77]
  assign _T_548 = _T_546[17:1]; // @[Shift.scala 90:30]
  assign _T_549 = _T_546[0:0]; // @[Shift.scala 90:48]
  assign _GEN_24 = {{16'd0}, _T_549}; // @[Shift.scala 90:39]
  assign _T_551 = _T_548 | _GEN_24; // @[Shift.scala 90:39]
  assign _T_553 = _T_546[17]; // @[Shift.scala 12:21]
  assign _T_554 = {_T_553,_T_551}; // @[Cat.scala 29:58]
  assign _T_555 = _T_547 ? _T_554 : _T_546; // @[Shift.scala 91:22]
  assign _T_558 = _T_509 ? 18'h3ffff : 18'h0; // @[Bitwise.scala 71:12]
  assign _T_559 = _T_502 ? _T_555 : _T_558; // @[Shift.scala 39:10]
  assign _T_560 = _T_559[3]; // @[convert.scala 55:31]
  assign _T_561 = _T_559[2]; // @[convert.scala 56:31]
  assign _T_562 = _T_559[1]; // @[convert.scala 57:31]
  assign _T_563 = _T_559[0]; // @[convert.scala 58:31]
  assign _T_564 = _T_559[17:3]; // @[convert.scala 59:69]
  assign _T_565 = _T_564 != 15'h0; // @[convert.scala 59:81]
  assign _T_566 = ~ _T_565; // @[convert.scala 59:50]
  assign _T_568 = _T_564 == 15'h7fff; // @[convert.scala 60:81]
  assign _T_569 = _T_560 | _T_562; // @[convert.scala 61:44]
  assign _T_570 = _T_569 | _T_563; // @[convert.scala 61:52]
  assign _T_571 = _T_561 & _T_570; // @[convert.scala 61:36]
  assign _T_572 = ~ _T_568; // @[convert.scala 62:63]
  assign _T_573 = _T_572 & _T_571; // @[convert.scala 62:103]
  assign _T_574 = _T_566 | _T_573; // @[convert.scala 62:60]
  assign _GEN_25 = {{14'd0}, _T_574}; // @[convert.scala 63:56]
  assign _T_577 = _T_564 + _GEN_25; // @[convert.scala 63:56]
  assign _T_578 = {decQ_sign,_T_577}; // @[Cat.scala 29:58]
  assign _T_580 = isZero_Z ? 16'h0 : _T_578; // @[Mux.scala 87:16]
  assign io_inReady = cycleNum <= 5'h1; // @[PositDivisionSqrt.scala 231:17]
  assign io_diviValid = outValid & _T_390; // @[PositDivisionSqrt.scala 232:17]
  assign io_sqrtValid = outValid & sqrtOp_Z; // @[PositDivisionSqrt.scala 233:17]
  assign io_invalidExc = isNaR_Z; // @[PositDivisionSqrt.scala 234:17]
  assign io_Q = isNaR_Z ? 16'h8000 : _T_580; // @[PositDivisionSqrt.scala 235:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleNum = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sqrtOp_Z = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  isNaR_Z = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  isZero_Z = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  scale_Z = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  signB_Z = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fractB_Z = _RAND_6[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rem_Z = _RAND_7[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sigX_Z = _RAND_8[18:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      cycleNum <= 5'h0;
    end else begin
      if (_T_349) begin
        cycleNum <= _T_366;
      end
    end
    if (entering) begin
      sqrtOp_Z <= io_sqrtOp;
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isNaR_Z <= _T_333;
      end else begin
        isNaR_Z <= _T_335;
      end
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isZero_Z <= decA_isZero;
      end else begin
        isZero_Z <= _T_339;
      end
    end
    if (entering_normalCase) begin
      if (io_sqrtOp) begin
        scale_Z <= {{2{_T_367[4]}},_T_367};
      end else begin
        scale_Z <= sExpQuot_S_div;
      end
    end
    if (_T_370) begin
      signB_Z <= _T_163;
    end
    if (_T_370) begin
      fractB_Z <= decB_fraction;
    end
    if (_T_443) begin
      if (ready) begin
        if (_T_410) begin
          rem_Z <= _T_413;
        end else begin
          rem_Z <= _T_415;
        end
      end else begin
        if (_T_410) begin
          rem_Z <= _T_424;
        end else begin
          rem_Z <= _T_428;
        end
      end
    end
    if (_T_447) begin
      sigX_Z <= _T_458;
    end
  end
endmodule
