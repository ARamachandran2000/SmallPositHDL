module PositAdder14_1(
  input         clock,
  input         reset,
  input  [13:0] io_A,
  input  [13:0] io_B,
  output [13:0] io_S
);
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [11:0] _T_4; // @[convert.scala 19:24]
  wire [11:0] _T_5; // @[convert.scala 19:43]
  wire [11:0] _T_6; // @[convert.scala 19:39]
  wire [7:0] _T_7; // @[LZD.scala 43:32]
  wire [3:0] _T_8; // @[LZD.scala 43:32]
  wire [1:0] _T_9; // @[LZD.scala 43:32]
  wire  _T_10; // @[LZD.scala 39:14]
  wire  _T_11; // @[LZD.scala 39:21]
  wire  _T_12; // @[LZD.scala 39:30]
  wire  _T_13; // @[LZD.scala 39:27]
  wire  _T_14; // @[LZD.scala 39:25]
  wire [1:0] _T_15; // @[Cat.scala 29:58]
  wire [1:0] _T_16; // @[LZD.scala 44:32]
  wire  _T_17; // @[LZD.scala 39:14]
  wire  _T_18; // @[LZD.scala 39:21]
  wire  _T_19; // @[LZD.scala 39:30]
  wire  _T_20; // @[LZD.scala 39:27]
  wire  _T_21; // @[LZD.scala 39:25]
  wire [1:0] _T_22; // @[Cat.scala 29:58]
  wire  _T_23; // @[Shift.scala 12:21]
  wire  _T_24; // @[Shift.scala 12:21]
  wire  _T_25; // @[LZD.scala 49:16]
  wire  _T_26; // @[LZD.scala 49:27]
  wire  _T_27; // @[LZD.scala 49:25]
  wire  _T_28; // @[LZD.scala 49:47]
  wire  _T_29; // @[LZD.scala 49:59]
  wire  _T_30; // @[LZD.scala 49:35]
  wire [2:0] _T_32; // @[Cat.scala 29:58]
  wire [3:0] _T_33; // @[LZD.scala 44:32]
  wire [1:0] _T_34; // @[LZD.scala 43:32]
  wire  _T_35; // @[LZD.scala 39:14]
  wire  _T_36; // @[LZD.scala 39:21]
  wire  _T_37; // @[LZD.scala 39:30]
  wire  _T_38; // @[LZD.scala 39:27]
  wire  _T_39; // @[LZD.scala 39:25]
  wire [1:0] _T_40; // @[Cat.scala 29:58]
  wire [1:0] _T_41; // @[LZD.scala 44:32]
  wire  _T_42; // @[LZD.scala 39:14]
  wire  _T_43; // @[LZD.scala 39:21]
  wire  _T_44; // @[LZD.scala 39:30]
  wire  _T_45; // @[LZD.scala 39:27]
  wire  _T_46; // @[LZD.scala 39:25]
  wire [1:0] _T_47; // @[Cat.scala 29:58]
  wire  _T_48; // @[Shift.scala 12:21]
  wire  _T_49; // @[Shift.scala 12:21]
  wire  _T_50; // @[LZD.scala 49:16]
  wire  _T_51; // @[LZD.scala 49:27]
  wire  _T_52; // @[LZD.scala 49:25]
  wire  _T_53; // @[LZD.scala 49:47]
  wire  _T_54; // @[LZD.scala 49:59]
  wire  _T_55; // @[LZD.scala 49:35]
  wire [2:0] _T_57; // @[Cat.scala 29:58]
  wire  _T_58; // @[Shift.scala 12:21]
  wire  _T_59; // @[Shift.scala 12:21]
  wire  _T_60; // @[LZD.scala 49:16]
  wire  _T_61; // @[LZD.scala 49:27]
  wire  _T_62; // @[LZD.scala 49:25]
  wire [1:0] _T_63; // @[LZD.scala 49:47]
  wire [1:0] _T_64; // @[LZD.scala 49:59]
  wire [1:0] _T_65; // @[LZD.scala 49:35]
  wire [3:0] _T_67; // @[Cat.scala 29:58]
  wire [3:0] _T_68; // @[LZD.scala 44:32]
  wire [1:0] _T_69; // @[LZD.scala 43:32]
  wire  _T_70; // @[LZD.scala 39:14]
  wire  _T_71; // @[LZD.scala 39:21]
  wire  _T_72; // @[LZD.scala 39:30]
  wire  _T_73; // @[LZD.scala 39:27]
  wire  _T_74; // @[LZD.scala 39:25]
  wire [1:0] _T_75; // @[Cat.scala 29:58]
  wire [1:0] _T_76; // @[LZD.scala 44:32]
  wire  _T_77; // @[LZD.scala 39:14]
  wire  _T_78; // @[LZD.scala 39:21]
  wire  _T_79; // @[LZD.scala 39:30]
  wire  _T_80; // @[LZD.scala 39:27]
  wire  _T_81; // @[LZD.scala 39:25]
  wire [1:0] _T_82; // @[Cat.scala 29:58]
  wire  _T_83; // @[Shift.scala 12:21]
  wire  _T_84; // @[Shift.scala 12:21]
  wire  _T_85; // @[LZD.scala 49:16]
  wire  _T_86; // @[LZD.scala 49:27]
  wire  _T_87; // @[LZD.scala 49:25]
  wire  _T_88; // @[LZD.scala 49:47]
  wire  _T_89; // @[LZD.scala 49:59]
  wire  _T_90; // @[LZD.scala 49:35]
  wire [2:0] _T_92; // @[Cat.scala 29:58]
  wire  _T_93; // @[Shift.scala 12:21]
  wire [2:0] _T_95; // @[LZD.scala 55:32]
  wire [2:0] _T_96; // @[LZD.scala 55:20]
  wire [3:0] _T_97; // @[Cat.scala 29:58]
  wire [3:0] _T_98; // @[convert.scala 21:22]
  wire [10:0] _T_99; // @[convert.scala 22:36]
  wire  _T_100; // @[Shift.scala 16:24]
  wire  _T_102; // @[Shift.scala 12:21]
  wire [2:0] _T_103; // @[Shift.scala 64:52]
  wire [10:0] _T_105; // @[Cat.scala 29:58]
  wire [10:0] _T_106; // @[Shift.scala 64:27]
  wire [2:0] _T_107; // @[Shift.scala 66:70]
  wire  _T_108; // @[Shift.scala 12:21]
  wire [6:0] _T_109; // @[Shift.scala 64:52]
  wire [10:0] _T_111; // @[Cat.scala 29:58]
  wire [10:0] _T_112; // @[Shift.scala 64:27]
  wire [1:0] _T_113; // @[Shift.scala 66:70]
  wire  _T_114; // @[Shift.scala 12:21]
  wire [8:0] _T_115; // @[Shift.scala 64:52]
  wire [10:0] _T_117; // @[Cat.scala 29:58]
  wire [10:0] _T_118; // @[Shift.scala 64:27]
  wire  _T_119; // @[Shift.scala 66:70]
  wire [9:0] _T_121; // @[Shift.scala 64:52]
  wire [10:0] _T_122; // @[Cat.scala 29:58]
  wire [10:0] _T_123; // @[Shift.scala 64:27]
  wire [10:0] _T_124; // @[Shift.scala 16:10]
  wire  _T_125; // @[convert.scala 23:34]
  wire [9:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_127; // @[convert.scala 25:26]
  wire [3:0] _T_129; // @[convert.scala 25:42]
  wire  _T_132; // @[convert.scala 26:67]
  wire  _T_133; // @[convert.scala 26:51]
  wire [5:0] _T_134; // @[Cat.scala 29:58]
  wire [12:0] _T_136; // @[convert.scala 29:56]
  wire  _T_137; // @[convert.scala 29:60]
  wire  _T_138; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_141; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [5:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_150; // @[convert.scala 18:24]
  wire  _T_151; // @[convert.scala 18:40]
  wire  _T_152; // @[convert.scala 18:36]
  wire [11:0] _T_153; // @[convert.scala 19:24]
  wire [11:0] _T_154; // @[convert.scala 19:43]
  wire [11:0] _T_155; // @[convert.scala 19:39]
  wire [7:0] _T_156; // @[LZD.scala 43:32]
  wire [3:0] _T_157; // @[LZD.scala 43:32]
  wire [1:0] _T_158; // @[LZD.scala 43:32]
  wire  _T_159; // @[LZD.scala 39:14]
  wire  _T_160; // @[LZD.scala 39:21]
  wire  _T_161; // @[LZD.scala 39:30]
  wire  _T_162; // @[LZD.scala 39:27]
  wire  _T_163; // @[LZD.scala 39:25]
  wire [1:0] _T_164; // @[Cat.scala 29:58]
  wire [1:0] _T_165; // @[LZD.scala 44:32]
  wire  _T_166; // @[LZD.scala 39:14]
  wire  _T_167; // @[LZD.scala 39:21]
  wire  _T_168; // @[LZD.scala 39:30]
  wire  _T_169; // @[LZD.scala 39:27]
  wire  _T_170; // @[LZD.scala 39:25]
  wire [1:0] _T_171; // @[Cat.scala 29:58]
  wire  _T_172; // @[Shift.scala 12:21]
  wire  _T_173; // @[Shift.scala 12:21]
  wire  _T_174; // @[LZD.scala 49:16]
  wire  _T_175; // @[LZD.scala 49:27]
  wire  _T_176; // @[LZD.scala 49:25]
  wire  _T_177; // @[LZD.scala 49:47]
  wire  _T_178; // @[LZD.scala 49:59]
  wire  _T_179; // @[LZD.scala 49:35]
  wire [2:0] _T_181; // @[Cat.scala 29:58]
  wire [3:0] _T_182; // @[LZD.scala 44:32]
  wire [1:0] _T_183; // @[LZD.scala 43:32]
  wire  _T_184; // @[LZD.scala 39:14]
  wire  _T_185; // @[LZD.scala 39:21]
  wire  _T_186; // @[LZD.scala 39:30]
  wire  _T_187; // @[LZD.scala 39:27]
  wire  _T_188; // @[LZD.scala 39:25]
  wire [1:0] _T_189; // @[Cat.scala 29:58]
  wire [1:0] _T_190; // @[LZD.scala 44:32]
  wire  _T_191; // @[LZD.scala 39:14]
  wire  _T_192; // @[LZD.scala 39:21]
  wire  _T_193; // @[LZD.scala 39:30]
  wire  _T_194; // @[LZD.scala 39:27]
  wire  _T_195; // @[LZD.scala 39:25]
  wire [1:0] _T_196; // @[Cat.scala 29:58]
  wire  _T_197; // @[Shift.scala 12:21]
  wire  _T_198; // @[Shift.scala 12:21]
  wire  _T_199; // @[LZD.scala 49:16]
  wire  _T_200; // @[LZD.scala 49:27]
  wire  _T_201; // @[LZD.scala 49:25]
  wire  _T_202; // @[LZD.scala 49:47]
  wire  _T_203; // @[LZD.scala 49:59]
  wire  _T_204; // @[LZD.scala 49:35]
  wire [2:0] _T_206; // @[Cat.scala 29:58]
  wire  _T_207; // @[Shift.scala 12:21]
  wire  _T_208; // @[Shift.scala 12:21]
  wire  _T_209; // @[LZD.scala 49:16]
  wire  _T_210; // @[LZD.scala 49:27]
  wire  _T_211; // @[LZD.scala 49:25]
  wire [1:0] _T_212; // @[LZD.scala 49:47]
  wire [1:0] _T_213; // @[LZD.scala 49:59]
  wire [1:0] _T_214; // @[LZD.scala 49:35]
  wire [3:0] _T_216; // @[Cat.scala 29:58]
  wire [3:0] _T_217; // @[LZD.scala 44:32]
  wire [1:0] _T_218; // @[LZD.scala 43:32]
  wire  _T_219; // @[LZD.scala 39:14]
  wire  _T_220; // @[LZD.scala 39:21]
  wire  _T_221; // @[LZD.scala 39:30]
  wire  _T_222; // @[LZD.scala 39:27]
  wire  _T_223; // @[LZD.scala 39:25]
  wire [1:0] _T_224; // @[Cat.scala 29:58]
  wire [1:0] _T_225; // @[LZD.scala 44:32]
  wire  _T_226; // @[LZD.scala 39:14]
  wire  _T_227; // @[LZD.scala 39:21]
  wire  _T_228; // @[LZD.scala 39:30]
  wire  _T_229; // @[LZD.scala 39:27]
  wire  _T_230; // @[LZD.scala 39:25]
  wire [1:0] _T_231; // @[Cat.scala 29:58]
  wire  _T_232; // @[Shift.scala 12:21]
  wire  _T_233; // @[Shift.scala 12:21]
  wire  _T_234; // @[LZD.scala 49:16]
  wire  _T_235; // @[LZD.scala 49:27]
  wire  _T_236; // @[LZD.scala 49:25]
  wire  _T_237; // @[LZD.scala 49:47]
  wire  _T_238; // @[LZD.scala 49:59]
  wire  _T_239; // @[LZD.scala 49:35]
  wire [2:0] _T_241; // @[Cat.scala 29:58]
  wire  _T_242; // @[Shift.scala 12:21]
  wire [2:0] _T_244; // @[LZD.scala 55:32]
  wire [2:0] _T_245; // @[LZD.scala 55:20]
  wire [3:0] _T_246; // @[Cat.scala 29:58]
  wire [3:0] _T_247; // @[convert.scala 21:22]
  wire [10:0] _T_248; // @[convert.scala 22:36]
  wire  _T_249; // @[Shift.scala 16:24]
  wire  _T_251; // @[Shift.scala 12:21]
  wire [2:0] _T_252; // @[Shift.scala 64:52]
  wire [10:0] _T_254; // @[Cat.scala 29:58]
  wire [10:0] _T_255; // @[Shift.scala 64:27]
  wire [2:0] _T_256; // @[Shift.scala 66:70]
  wire  _T_257; // @[Shift.scala 12:21]
  wire [6:0] _T_258; // @[Shift.scala 64:52]
  wire [10:0] _T_260; // @[Cat.scala 29:58]
  wire [10:0] _T_261; // @[Shift.scala 64:27]
  wire [1:0] _T_262; // @[Shift.scala 66:70]
  wire  _T_263; // @[Shift.scala 12:21]
  wire [8:0] _T_264; // @[Shift.scala 64:52]
  wire [10:0] _T_266; // @[Cat.scala 29:58]
  wire [10:0] _T_267; // @[Shift.scala 64:27]
  wire  _T_268; // @[Shift.scala 66:70]
  wire [9:0] _T_270; // @[Shift.scala 64:52]
  wire [10:0] _T_271; // @[Cat.scala 29:58]
  wire [10:0] _T_272; // @[Shift.scala 64:27]
  wire [10:0] _T_273; // @[Shift.scala 16:10]
  wire  _T_274; // @[convert.scala 23:34]
  wire [9:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_276; // @[convert.scala 25:26]
  wire [3:0] _T_278; // @[convert.scala 25:42]
  wire  _T_281; // @[convert.scala 26:67]
  wire  _T_282; // @[convert.scala 26:51]
  wire [5:0] _T_283; // @[Cat.scala 29:58]
  wire [12:0] _T_285; // @[convert.scala 29:56]
  wire  _T_286; // @[convert.scala 29:60]
  wire  _T_287; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_290; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [5:0] decB_scale; // @[convert.scala 32:24]
  wire  aGTb; // @[PositAdder.scala 24:32]
  wire  greaterSign; // @[PositAdder.scala 25:24]
  wire  smallerSign; // @[PositAdder.scala 26:24]
  wire [5:0] greaterExp; // @[PositAdder.scala 27:24]
  wire [5:0] smallerExp; // @[PositAdder.scala 28:24]
  wire [9:0] greaterFrac; // @[PositAdder.scala 29:24]
  wire [9:0] smallerFrac; // @[PositAdder.scala 30:24]
  wire  smallerZero; // @[PositAdder.scala 31:24]
  wire [5:0] _T_299; // @[PositAdder.scala 32:32]
  wire [5:0] scale_diff; // @[PositAdder.scala 32:32]
  wire  _T_300; // @[PositAdder.scala 33:38]
  wire [11:0] greaterSig; // @[Cat.scala 29:58]
  wire  _T_302; // @[PositAdder.scala 34:52]
  wire  _T_303; // @[PositAdder.scala 34:38]
  wire [14:0] _T_306; // @[Cat.scala 29:58]
  wire [5:0] _T_307; // @[PositAdder.scala 35:68]
  wire  _T_308; // @[Shift.scala 39:24]
  wire [3:0] _T_309; // @[Shift.scala 40:44]
  wire [6:0] _T_310; // @[Shift.scala 90:30]
  wire [7:0] _T_311; // @[Shift.scala 90:48]
  wire  _T_312; // @[Shift.scala 90:57]
  wire [6:0] _GEN_0; // @[Shift.scala 90:39]
  wire [6:0] _T_313; // @[Shift.scala 90:39]
  wire  _T_314; // @[Shift.scala 12:21]
  wire  _T_315; // @[Shift.scala 12:21]
  wire [7:0] _T_317; // @[Bitwise.scala 71:12]
  wire [14:0] _T_318; // @[Cat.scala 29:58]
  wire [14:0] _T_319; // @[Shift.scala 91:22]
  wire [2:0] _T_320; // @[Shift.scala 92:77]
  wire [10:0] _T_321; // @[Shift.scala 90:30]
  wire [3:0] _T_322; // @[Shift.scala 90:48]
  wire  _T_323; // @[Shift.scala 90:57]
  wire [10:0] _GEN_1; // @[Shift.scala 90:39]
  wire [10:0] _T_324; // @[Shift.scala 90:39]
  wire  _T_325; // @[Shift.scala 12:21]
  wire  _T_326; // @[Shift.scala 12:21]
  wire [3:0] _T_328; // @[Bitwise.scala 71:12]
  wire [14:0] _T_329; // @[Cat.scala 29:58]
  wire [14:0] _T_330; // @[Shift.scala 91:22]
  wire [1:0] _T_331; // @[Shift.scala 92:77]
  wire [12:0] _T_332; // @[Shift.scala 90:30]
  wire [1:0] _T_333; // @[Shift.scala 90:48]
  wire  _T_334; // @[Shift.scala 90:57]
  wire [12:0] _GEN_2; // @[Shift.scala 90:39]
  wire [12:0] _T_335; // @[Shift.scala 90:39]
  wire  _T_336; // @[Shift.scala 12:21]
  wire  _T_337; // @[Shift.scala 12:21]
  wire [1:0] _T_339; // @[Bitwise.scala 71:12]
  wire [14:0] _T_340; // @[Cat.scala 29:58]
  wire [14:0] _T_341; // @[Shift.scala 91:22]
  wire  _T_342; // @[Shift.scala 92:77]
  wire [13:0] _T_343; // @[Shift.scala 90:30]
  wire  _T_344; // @[Shift.scala 90:48]
  wire [13:0] _GEN_3; // @[Shift.scala 90:39]
  wire [13:0] _T_346; // @[Shift.scala 90:39]
  wire  _T_348; // @[Shift.scala 12:21]
  wire [14:0] _T_349; // @[Cat.scala 29:58]
  wire [14:0] _T_350; // @[Shift.scala 91:22]
  wire [14:0] _T_353; // @[Bitwise.scala 71:12]
  wire [14:0] smallerSig; // @[Shift.scala 39:10]
  wire [11:0] _T_354; // @[PositAdder.scala 36:45]
  wire [12:0] rawSumSig; // @[PositAdder.scala 36:32]
  wire  _T_355; // @[PositAdder.scala 37:31]
  wire  _T_356; // @[PositAdder.scala 37:59]
  wire  sumSign; // @[PositAdder.scala 37:43]
  wire [11:0] _T_357; // @[PositAdder.scala 38:48]
  wire [2:0] _T_358; // @[PositAdder.scala 38:63]
  wire [15:0] signSumSig; // @[Cat.scala 29:58]
  wire [14:0] _T_360; // @[PositAdder.scala 40:31]
  wire [14:0] _T_361; // @[PositAdder.scala 40:66]
  wire [14:0] sumXor; // @[PositAdder.scala 40:49]
  wire [7:0] _T_362; // @[LZD.scala 43:32]
  wire [3:0] _T_363; // @[LZD.scala 43:32]
  wire [1:0] _T_364; // @[LZD.scala 43:32]
  wire  _T_365; // @[LZD.scala 39:14]
  wire  _T_366; // @[LZD.scala 39:21]
  wire  _T_367; // @[LZD.scala 39:30]
  wire  _T_368; // @[LZD.scala 39:27]
  wire  _T_369; // @[LZD.scala 39:25]
  wire [1:0] _T_370; // @[Cat.scala 29:58]
  wire [1:0] _T_371; // @[LZD.scala 44:32]
  wire  _T_372; // @[LZD.scala 39:14]
  wire  _T_373; // @[LZD.scala 39:21]
  wire  _T_374; // @[LZD.scala 39:30]
  wire  _T_375; // @[LZD.scala 39:27]
  wire  _T_376; // @[LZD.scala 39:25]
  wire [1:0] _T_377; // @[Cat.scala 29:58]
  wire  _T_378; // @[Shift.scala 12:21]
  wire  _T_379; // @[Shift.scala 12:21]
  wire  _T_380; // @[LZD.scala 49:16]
  wire  _T_381; // @[LZD.scala 49:27]
  wire  _T_382; // @[LZD.scala 49:25]
  wire  _T_383; // @[LZD.scala 49:47]
  wire  _T_384; // @[LZD.scala 49:59]
  wire  _T_385; // @[LZD.scala 49:35]
  wire [2:0] _T_387; // @[Cat.scala 29:58]
  wire [3:0] _T_388; // @[LZD.scala 44:32]
  wire [1:0] _T_389; // @[LZD.scala 43:32]
  wire  _T_390; // @[LZD.scala 39:14]
  wire  _T_391; // @[LZD.scala 39:21]
  wire  _T_392; // @[LZD.scala 39:30]
  wire  _T_393; // @[LZD.scala 39:27]
  wire  _T_394; // @[LZD.scala 39:25]
  wire [1:0] _T_395; // @[Cat.scala 29:58]
  wire [1:0] _T_396; // @[LZD.scala 44:32]
  wire  _T_397; // @[LZD.scala 39:14]
  wire  _T_398; // @[LZD.scala 39:21]
  wire  _T_399; // @[LZD.scala 39:30]
  wire  _T_400; // @[LZD.scala 39:27]
  wire  _T_401; // @[LZD.scala 39:25]
  wire [1:0] _T_402; // @[Cat.scala 29:58]
  wire  _T_403; // @[Shift.scala 12:21]
  wire  _T_404; // @[Shift.scala 12:21]
  wire  _T_405; // @[LZD.scala 49:16]
  wire  _T_406; // @[LZD.scala 49:27]
  wire  _T_407; // @[LZD.scala 49:25]
  wire  _T_408; // @[LZD.scala 49:47]
  wire  _T_409; // @[LZD.scala 49:59]
  wire  _T_410; // @[LZD.scala 49:35]
  wire [2:0] _T_412; // @[Cat.scala 29:58]
  wire  _T_413; // @[Shift.scala 12:21]
  wire  _T_414; // @[Shift.scala 12:21]
  wire  _T_415; // @[LZD.scala 49:16]
  wire  _T_416; // @[LZD.scala 49:27]
  wire  _T_417; // @[LZD.scala 49:25]
  wire [1:0] _T_418; // @[LZD.scala 49:47]
  wire [1:0] _T_419; // @[LZD.scala 49:59]
  wire [1:0] _T_420; // @[LZD.scala 49:35]
  wire [3:0] _T_422; // @[Cat.scala 29:58]
  wire [6:0] _T_423; // @[LZD.scala 44:32]
  wire [3:0] _T_424; // @[LZD.scala 43:32]
  wire [1:0] _T_425; // @[LZD.scala 43:32]
  wire  _T_426; // @[LZD.scala 39:14]
  wire  _T_427; // @[LZD.scala 39:21]
  wire  _T_428; // @[LZD.scala 39:30]
  wire  _T_429; // @[LZD.scala 39:27]
  wire  _T_430; // @[LZD.scala 39:25]
  wire [1:0] _T_431; // @[Cat.scala 29:58]
  wire [1:0] _T_432; // @[LZD.scala 44:32]
  wire  _T_433; // @[LZD.scala 39:14]
  wire  _T_434; // @[LZD.scala 39:21]
  wire  _T_435; // @[LZD.scala 39:30]
  wire  _T_436; // @[LZD.scala 39:27]
  wire  _T_437; // @[LZD.scala 39:25]
  wire [1:0] _T_438; // @[Cat.scala 29:58]
  wire  _T_439; // @[Shift.scala 12:21]
  wire  _T_440; // @[Shift.scala 12:21]
  wire  _T_441; // @[LZD.scala 49:16]
  wire  _T_442; // @[LZD.scala 49:27]
  wire  _T_443; // @[LZD.scala 49:25]
  wire  _T_444; // @[LZD.scala 49:47]
  wire  _T_445; // @[LZD.scala 49:59]
  wire  _T_446; // @[LZD.scala 49:35]
  wire [2:0] _T_448; // @[Cat.scala 29:58]
  wire [2:0] _T_449; // @[LZD.scala 44:32]
  wire [1:0] _T_450; // @[LZD.scala 43:32]
  wire  _T_451; // @[LZD.scala 39:14]
  wire  _T_452; // @[LZD.scala 39:21]
  wire  _T_453; // @[LZD.scala 39:30]
  wire  _T_454; // @[LZD.scala 39:27]
  wire  _T_455; // @[LZD.scala 39:25]
  wire [1:0] _T_456; // @[Cat.scala 29:58]
  wire  _T_457; // @[LZD.scala 44:32]
  wire  _T_459; // @[Shift.scala 12:21]
  wire  _T_461; // @[LZD.scala 55:32]
  wire  _T_462; // @[LZD.scala 55:20]
  wire [1:0] _T_463; // @[Cat.scala 29:58]
  wire  _T_464; // @[Shift.scala 12:21]
  wire [1:0] _T_466; // @[LZD.scala 55:32]
  wire [1:0] _T_467; // @[LZD.scala 55:20]
  wire [2:0] _T_468; // @[Cat.scala 29:58]
  wire  _T_469; // @[Shift.scala 12:21]
  wire [2:0] _T_471; // @[LZD.scala 55:32]
  wire [2:0] _T_472; // @[LZD.scala 55:20]
  wire [3:0] sumLZD; // @[Cat.scala 29:58]
  wire [4:0] _T_473; // @[Cat.scala 29:58]
  wire [4:0] _T_474; // @[PositAdder.scala 42:38]
  wire [4:0] _T_476; // @[PositAdder.scala 42:45]
  wire [4:0] scaleBias; // @[PositAdder.scala 42:45]
  wire [5:0] _GEN_4; // @[PositAdder.scala 43:32]
  wire [6:0] sumScale; // @[PositAdder.scala 43:32]
  wire  overflow; // @[PositAdder.scala 44:30]
  wire [3:0] normalShift; // @[PositAdder.scala 45:22]
  wire [13:0] _T_477; // @[PositAdder.scala 46:36]
  wire  _T_478; // @[Shift.scala 16:24]
  wire  _T_480; // @[Shift.scala 12:21]
  wire [5:0] _T_481; // @[Shift.scala 64:52]
  wire [13:0] _T_483; // @[Cat.scala 29:58]
  wire [13:0] _T_484; // @[Shift.scala 64:27]
  wire [2:0] _T_485; // @[Shift.scala 66:70]
  wire  _T_486; // @[Shift.scala 12:21]
  wire [9:0] _T_487; // @[Shift.scala 64:52]
  wire [13:0] _T_489; // @[Cat.scala 29:58]
  wire [13:0] _T_490; // @[Shift.scala 64:27]
  wire [1:0] _T_491; // @[Shift.scala 66:70]
  wire  _T_492; // @[Shift.scala 12:21]
  wire [11:0] _T_493; // @[Shift.scala 64:52]
  wire [13:0] _T_495; // @[Cat.scala 29:58]
  wire [13:0] _T_496; // @[Shift.scala 64:27]
  wire  _T_497; // @[Shift.scala 66:70]
  wire [12:0] _T_499; // @[Shift.scala 64:52]
  wire [13:0] _T_500; // @[Cat.scala 29:58]
  wire [13:0] _T_501; // @[Shift.scala 64:27]
  wire [13:0] shiftSig; // @[Shift.scala 16:10]
  wire [6:0] _T_502; // @[PositAdder.scala 51:24]
  wire [9:0] decS_fraction; // @[PositAdder.scala 52:34]
  wire  decS_isNaR; // @[PositAdder.scala 53:32]
  wire  _T_505; // @[PositAdder.scala 54:33]
  wire  _T_506; // @[PositAdder.scala 54:21]
  wire  _T_507; // @[PositAdder.scala 54:52]
  wire  decS_isZero; // @[PositAdder.scala 54:37]
  wire [1:0] _T_509; // @[PositAdder.scala 55:33]
  wire  _T_510; // @[PositAdder.scala 55:49]
  wire  _T_511; // @[PositAdder.scala 55:63]
  wire  _T_512; // @[PositAdder.scala 55:53]
  wire [5:0] _GEN_5; // @[PositAdder.scala 48:25 PositAdder.scala 51:18]
  wire [5:0] decS_scale; // @[PositAdder.scala 48:25 PositAdder.scala 51:18]
  wire  _T_515; // @[convert.scala 46:61]
  wire  _T_516; // @[convert.scala 46:52]
  wire  _T_518; // @[convert.scala 46:42]
  wire [4:0] _T_519; // @[convert.scala 48:34]
  wire  _T_520; // @[convert.scala 49:36]
  wire [4:0] _T_522; // @[convert.scala 50:36]
  wire [4:0] _T_523; // @[convert.scala 50:36]
  wire [4:0] _T_524; // @[convert.scala 50:28]
  wire  _T_525; // @[convert.scala 51:31]
  wire  _T_526; // @[convert.scala 52:43]
  wire [15:0] _T_530; // @[Cat.scala 29:58]
  wire [4:0] _T_531; // @[Shift.scala 39:17]
  wire  _T_532; // @[Shift.scala 39:24]
  wire [3:0] _T_533; // @[Shift.scala 40:44]
  wire [7:0] _T_534; // @[Shift.scala 90:30]
  wire [7:0] _T_535; // @[Shift.scala 90:48]
  wire  _T_536; // @[Shift.scala 90:57]
  wire [7:0] _GEN_6; // @[Shift.scala 90:39]
  wire [7:0] _T_537; // @[Shift.scala 90:39]
  wire  _T_538; // @[Shift.scala 12:21]
  wire  _T_539; // @[Shift.scala 12:21]
  wire [7:0] _T_541; // @[Bitwise.scala 71:12]
  wire [15:0] _T_542; // @[Cat.scala 29:58]
  wire [15:0] _T_543; // @[Shift.scala 91:22]
  wire [2:0] _T_544; // @[Shift.scala 92:77]
  wire [11:0] _T_545; // @[Shift.scala 90:30]
  wire [3:0] _T_546; // @[Shift.scala 90:48]
  wire  _T_547; // @[Shift.scala 90:57]
  wire [11:0] _GEN_7; // @[Shift.scala 90:39]
  wire [11:0] _T_548; // @[Shift.scala 90:39]
  wire  _T_549; // @[Shift.scala 12:21]
  wire  _T_550; // @[Shift.scala 12:21]
  wire [3:0] _T_552; // @[Bitwise.scala 71:12]
  wire [15:0] _T_553; // @[Cat.scala 29:58]
  wire [15:0] _T_554; // @[Shift.scala 91:22]
  wire [1:0] _T_555; // @[Shift.scala 92:77]
  wire [13:0] _T_556; // @[Shift.scala 90:30]
  wire [1:0] _T_557; // @[Shift.scala 90:48]
  wire  _T_558; // @[Shift.scala 90:57]
  wire [13:0] _GEN_8; // @[Shift.scala 90:39]
  wire [13:0] _T_559; // @[Shift.scala 90:39]
  wire  _T_560; // @[Shift.scala 12:21]
  wire  _T_561; // @[Shift.scala 12:21]
  wire [1:0] _T_563; // @[Bitwise.scala 71:12]
  wire [15:0] _T_564; // @[Cat.scala 29:58]
  wire [15:0] _T_565; // @[Shift.scala 91:22]
  wire  _T_566; // @[Shift.scala 92:77]
  wire [14:0] _T_567; // @[Shift.scala 90:30]
  wire  _T_568; // @[Shift.scala 90:48]
  wire [14:0] _GEN_9; // @[Shift.scala 90:39]
  wire [14:0] _T_570; // @[Shift.scala 90:39]
  wire  _T_572; // @[Shift.scala 12:21]
  wire [15:0] _T_573; // @[Cat.scala 29:58]
  wire [15:0] _T_574; // @[Shift.scala 91:22]
  wire [15:0] _T_577; // @[Bitwise.scala 71:12]
  wire [15:0] _T_578; // @[Shift.scala 39:10]
  wire  _T_579; // @[convert.scala 55:31]
  wire  _T_580; // @[convert.scala 56:31]
  wire  _T_581; // @[convert.scala 57:31]
  wire  _T_582; // @[convert.scala 58:31]
  wire [12:0] _T_583; // @[convert.scala 59:69]
  wire  _T_584; // @[convert.scala 59:81]
  wire  _T_585; // @[convert.scala 59:50]
  wire  _T_587; // @[convert.scala 60:81]
  wire  _T_588; // @[convert.scala 61:44]
  wire  _T_589; // @[convert.scala 61:52]
  wire  _T_590; // @[convert.scala 61:36]
  wire  _T_591; // @[convert.scala 62:63]
  wire  _T_592; // @[convert.scala 62:103]
  wire  _T_593; // @[convert.scala 62:60]
  wire [12:0] _GEN_10; // @[convert.scala 63:56]
  wire [12:0] _T_596; // @[convert.scala 63:56]
  wire [13:0] _T_597; // @[Cat.scala 29:58]
  wire [13:0] _T_599; // @[Mux.scala 87:16]
  assign _T_1 = io_A[13]; // @[convert.scala 18:24]
  assign _T_2 = io_A[12]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[12:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[11:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[11:4]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[7:4]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8[3:2]; // @[LZD.scala 43:32]
  assign _T_10 = _T_9 != 2'h0; // @[LZD.scala 39:14]
  assign _T_11 = _T_9[1]; // @[LZD.scala 39:21]
  assign _T_12 = _T_9[0]; // @[LZD.scala 39:30]
  assign _T_13 = ~ _T_12; // @[LZD.scala 39:27]
  assign _T_14 = _T_11 | _T_13; // @[LZD.scala 39:25]
  assign _T_15 = {_T_10,_T_14}; // @[Cat.scala 29:58]
  assign _T_16 = _T_8[1:0]; // @[LZD.scala 44:32]
  assign _T_17 = _T_16 != 2'h0; // @[LZD.scala 39:14]
  assign _T_18 = _T_16[1]; // @[LZD.scala 39:21]
  assign _T_19 = _T_16[0]; // @[LZD.scala 39:30]
  assign _T_20 = ~ _T_19; // @[LZD.scala 39:27]
  assign _T_21 = _T_18 | _T_20; // @[LZD.scala 39:25]
  assign _T_22 = {_T_17,_T_21}; // @[Cat.scala 29:58]
  assign _T_23 = _T_15[1]; // @[Shift.scala 12:21]
  assign _T_24 = _T_22[1]; // @[Shift.scala 12:21]
  assign _T_25 = _T_23 | _T_24; // @[LZD.scala 49:16]
  assign _T_26 = ~ _T_24; // @[LZD.scala 49:27]
  assign _T_27 = _T_23 | _T_26; // @[LZD.scala 49:25]
  assign _T_28 = _T_15[0:0]; // @[LZD.scala 49:47]
  assign _T_29 = _T_22[0:0]; // @[LZD.scala 49:59]
  assign _T_30 = _T_23 ? _T_28 : _T_29; // @[LZD.scala 49:35]
  assign _T_32 = {_T_25,_T_27,_T_30}; // @[Cat.scala 29:58]
  assign _T_33 = _T_7[3:0]; // @[LZD.scala 44:32]
  assign _T_34 = _T_33[3:2]; // @[LZD.scala 43:32]
  assign _T_35 = _T_34 != 2'h0; // @[LZD.scala 39:14]
  assign _T_36 = _T_34[1]; // @[LZD.scala 39:21]
  assign _T_37 = _T_34[0]; // @[LZD.scala 39:30]
  assign _T_38 = ~ _T_37; // @[LZD.scala 39:27]
  assign _T_39 = _T_36 | _T_38; // @[LZD.scala 39:25]
  assign _T_40 = {_T_35,_T_39}; // @[Cat.scala 29:58]
  assign _T_41 = _T_33[1:0]; // @[LZD.scala 44:32]
  assign _T_42 = _T_41 != 2'h0; // @[LZD.scala 39:14]
  assign _T_43 = _T_41[1]; // @[LZD.scala 39:21]
  assign _T_44 = _T_41[0]; // @[LZD.scala 39:30]
  assign _T_45 = ~ _T_44; // @[LZD.scala 39:27]
  assign _T_46 = _T_43 | _T_45; // @[LZD.scala 39:25]
  assign _T_47 = {_T_42,_T_46}; // @[Cat.scala 29:58]
  assign _T_48 = _T_40[1]; // @[Shift.scala 12:21]
  assign _T_49 = _T_47[1]; // @[Shift.scala 12:21]
  assign _T_50 = _T_48 | _T_49; // @[LZD.scala 49:16]
  assign _T_51 = ~ _T_49; // @[LZD.scala 49:27]
  assign _T_52 = _T_48 | _T_51; // @[LZD.scala 49:25]
  assign _T_53 = _T_40[0:0]; // @[LZD.scala 49:47]
  assign _T_54 = _T_47[0:0]; // @[LZD.scala 49:59]
  assign _T_55 = _T_48 ? _T_53 : _T_54; // @[LZD.scala 49:35]
  assign _T_57 = {_T_50,_T_52,_T_55}; // @[Cat.scala 29:58]
  assign _T_58 = _T_32[2]; // @[Shift.scala 12:21]
  assign _T_59 = _T_57[2]; // @[Shift.scala 12:21]
  assign _T_60 = _T_58 | _T_59; // @[LZD.scala 49:16]
  assign _T_61 = ~ _T_59; // @[LZD.scala 49:27]
  assign _T_62 = _T_58 | _T_61; // @[LZD.scala 49:25]
  assign _T_63 = _T_32[1:0]; // @[LZD.scala 49:47]
  assign _T_64 = _T_57[1:0]; // @[LZD.scala 49:59]
  assign _T_65 = _T_58 ? _T_63 : _T_64; // @[LZD.scala 49:35]
  assign _T_67 = {_T_60,_T_62,_T_65}; // @[Cat.scala 29:58]
  assign _T_68 = _T_6[3:0]; // @[LZD.scala 44:32]
  assign _T_69 = _T_68[3:2]; // @[LZD.scala 43:32]
  assign _T_70 = _T_69 != 2'h0; // @[LZD.scala 39:14]
  assign _T_71 = _T_69[1]; // @[LZD.scala 39:21]
  assign _T_72 = _T_69[0]; // @[LZD.scala 39:30]
  assign _T_73 = ~ _T_72; // @[LZD.scala 39:27]
  assign _T_74 = _T_71 | _T_73; // @[LZD.scala 39:25]
  assign _T_75 = {_T_70,_T_74}; // @[Cat.scala 29:58]
  assign _T_76 = _T_68[1:0]; // @[LZD.scala 44:32]
  assign _T_77 = _T_76 != 2'h0; // @[LZD.scala 39:14]
  assign _T_78 = _T_76[1]; // @[LZD.scala 39:21]
  assign _T_79 = _T_76[0]; // @[LZD.scala 39:30]
  assign _T_80 = ~ _T_79; // @[LZD.scala 39:27]
  assign _T_81 = _T_78 | _T_80; // @[LZD.scala 39:25]
  assign _T_82 = {_T_77,_T_81}; // @[Cat.scala 29:58]
  assign _T_83 = _T_75[1]; // @[Shift.scala 12:21]
  assign _T_84 = _T_82[1]; // @[Shift.scala 12:21]
  assign _T_85 = _T_83 | _T_84; // @[LZD.scala 49:16]
  assign _T_86 = ~ _T_84; // @[LZD.scala 49:27]
  assign _T_87 = _T_83 | _T_86; // @[LZD.scala 49:25]
  assign _T_88 = _T_75[0:0]; // @[LZD.scala 49:47]
  assign _T_89 = _T_82[0:0]; // @[LZD.scala 49:59]
  assign _T_90 = _T_83 ? _T_88 : _T_89; // @[LZD.scala 49:35]
  assign _T_92 = {_T_85,_T_87,_T_90}; // @[Cat.scala 29:58]
  assign _T_93 = _T_67[3]; // @[Shift.scala 12:21]
  assign _T_95 = _T_67[2:0]; // @[LZD.scala 55:32]
  assign _T_96 = _T_93 ? _T_95 : _T_92; // @[LZD.scala 55:20]
  assign _T_97 = {_T_93,_T_96}; // @[Cat.scala 29:58]
  assign _T_98 = ~ _T_97; // @[convert.scala 21:22]
  assign _T_99 = io_A[10:0]; // @[convert.scala 22:36]
  assign _T_100 = _T_98 < 4'hb; // @[Shift.scala 16:24]
  assign _T_102 = _T_98[3]; // @[Shift.scala 12:21]
  assign _T_103 = _T_99[2:0]; // @[Shift.scala 64:52]
  assign _T_105 = {_T_103,8'h0}; // @[Cat.scala 29:58]
  assign _T_106 = _T_102 ? _T_105 : _T_99; // @[Shift.scala 64:27]
  assign _T_107 = _T_98[2:0]; // @[Shift.scala 66:70]
  assign _T_108 = _T_107[2]; // @[Shift.scala 12:21]
  assign _T_109 = _T_106[6:0]; // @[Shift.scala 64:52]
  assign _T_111 = {_T_109,4'h0}; // @[Cat.scala 29:58]
  assign _T_112 = _T_108 ? _T_111 : _T_106; // @[Shift.scala 64:27]
  assign _T_113 = _T_107[1:0]; // @[Shift.scala 66:70]
  assign _T_114 = _T_113[1]; // @[Shift.scala 12:21]
  assign _T_115 = _T_112[8:0]; // @[Shift.scala 64:52]
  assign _T_117 = {_T_115,2'h0}; // @[Cat.scala 29:58]
  assign _T_118 = _T_114 ? _T_117 : _T_112; // @[Shift.scala 64:27]
  assign _T_119 = _T_113[0:0]; // @[Shift.scala 66:70]
  assign _T_121 = _T_118[9:0]; // @[Shift.scala 64:52]
  assign _T_122 = {_T_121,1'h0}; // @[Cat.scala 29:58]
  assign _T_123 = _T_119 ? _T_122 : _T_118; // @[Shift.scala 64:27]
  assign _T_124 = _T_100 ? _T_123 : 11'h0; // @[Shift.scala 16:10]
  assign _T_125 = _T_124[10:10]; // @[convert.scala 23:34]
  assign decA_fraction = _T_124[9:0]; // @[convert.scala 24:34]
  assign _T_127 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_129 = _T_3 ? _T_98 : _T_97; // @[convert.scala 25:42]
  assign _T_132 = ~ _T_125; // @[convert.scala 26:67]
  assign _T_133 = _T_1 ? _T_132 : _T_125; // @[convert.scala 26:51]
  assign _T_134 = {_T_127,_T_129,_T_133}; // @[Cat.scala 29:58]
  assign _T_136 = io_A[12:0]; // @[convert.scala 29:56]
  assign _T_137 = _T_136 != 13'h0; // @[convert.scala 29:60]
  assign _T_138 = ~ _T_137; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_138; // @[convert.scala 29:39]
  assign _T_141 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_141 & _T_138; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_134); // @[convert.scala 32:24]
  assign _T_150 = io_B[13]; // @[convert.scala 18:24]
  assign _T_151 = io_B[12]; // @[convert.scala 18:40]
  assign _T_152 = _T_150 ^ _T_151; // @[convert.scala 18:36]
  assign _T_153 = io_B[12:1]; // @[convert.scala 19:24]
  assign _T_154 = io_B[11:0]; // @[convert.scala 19:43]
  assign _T_155 = _T_153 ^ _T_154; // @[convert.scala 19:39]
  assign _T_156 = _T_155[11:4]; // @[LZD.scala 43:32]
  assign _T_157 = _T_156[7:4]; // @[LZD.scala 43:32]
  assign _T_158 = _T_157[3:2]; // @[LZD.scala 43:32]
  assign _T_159 = _T_158 != 2'h0; // @[LZD.scala 39:14]
  assign _T_160 = _T_158[1]; // @[LZD.scala 39:21]
  assign _T_161 = _T_158[0]; // @[LZD.scala 39:30]
  assign _T_162 = ~ _T_161; // @[LZD.scala 39:27]
  assign _T_163 = _T_160 | _T_162; // @[LZD.scala 39:25]
  assign _T_164 = {_T_159,_T_163}; // @[Cat.scala 29:58]
  assign _T_165 = _T_157[1:0]; // @[LZD.scala 44:32]
  assign _T_166 = _T_165 != 2'h0; // @[LZD.scala 39:14]
  assign _T_167 = _T_165[1]; // @[LZD.scala 39:21]
  assign _T_168 = _T_165[0]; // @[LZD.scala 39:30]
  assign _T_169 = ~ _T_168; // @[LZD.scala 39:27]
  assign _T_170 = _T_167 | _T_169; // @[LZD.scala 39:25]
  assign _T_171 = {_T_166,_T_170}; // @[Cat.scala 29:58]
  assign _T_172 = _T_164[1]; // @[Shift.scala 12:21]
  assign _T_173 = _T_171[1]; // @[Shift.scala 12:21]
  assign _T_174 = _T_172 | _T_173; // @[LZD.scala 49:16]
  assign _T_175 = ~ _T_173; // @[LZD.scala 49:27]
  assign _T_176 = _T_172 | _T_175; // @[LZD.scala 49:25]
  assign _T_177 = _T_164[0:0]; // @[LZD.scala 49:47]
  assign _T_178 = _T_171[0:0]; // @[LZD.scala 49:59]
  assign _T_179 = _T_172 ? _T_177 : _T_178; // @[LZD.scala 49:35]
  assign _T_181 = {_T_174,_T_176,_T_179}; // @[Cat.scala 29:58]
  assign _T_182 = _T_156[3:0]; // @[LZD.scala 44:32]
  assign _T_183 = _T_182[3:2]; // @[LZD.scala 43:32]
  assign _T_184 = _T_183 != 2'h0; // @[LZD.scala 39:14]
  assign _T_185 = _T_183[1]; // @[LZD.scala 39:21]
  assign _T_186 = _T_183[0]; // @[LZD.scala 39:30]
  assign _T_187 = ~ _T_186; // @[LZD.scala 39:27]
  assign _T_188 = _T_185 | _T_187; // @[LZD.scala 39:25]
  assign _T_189 = {_T_184,_T_188}; // @[Cat.scala 29:58]
  assign _T_190 = _T_182[1:0]; // @[LZD.scala 44:32]
  assign _T_191 = _T_190 != 2'h0; // @[LZD.scala 39:14]
  assign _T_192 = _T_190[1]; // @[LZD.scala 39:21]
  assign _T_193 = _T_190[0]; // @[LZD.scala 39:30]
  assign _T_194 = ~ _T_193; // @[LZD.scala 39:27]
  assign _T_195 = _T_192 | _T_194; // @[LZD.scala 39:25]
  assign _T_196 = {_T_191,_T_195}; // @[Cat.scala 29:58]
  assign _T_197 = _T_189[1]; // @[Shift.scala 12:21]
  assign _T_198 = _T_196[1]; // @[Shift.scala 12:21]
  assign _T_199 = _T_197 | _T_198; // @[LZD.scala 49:16]
  assign _T_200 = ~ _T_198; // @[LZD.scala 49:27]
  assign _T_201 = _T_197 | _T_200; // @[LZD.scala 49:25]
  assign _T_202 = _T_189[0:0]; // @[LZD.scala 49:47]
  assign _T_203 = _T_196[0:0]; // @[LZD.scala 49:59]
  assign _T_204 = _T_197 ? _T_202 : _T_203; // @[LZD.scala 49:35]
  assign _T_206 = {_T_199,_T_201,_T_204}; // @[Cat.scala 29:58]
  assign _T_207 = _T_181[2]; // @[Shift.scala 12:21]
  assign _T_208 = _T_206[2]; // @[Shift.scala 12:21]
  assign _T_209 = _T_207 | _T_208; // @[LZD.scala 49:16]
  assign _T_210 = ~ _T_208; // @[LZD.scala 49:27]
  assign _T_211 = _T_207 | _T_210; // @[LZD.scala 49:25]
  assign _T_212 = _T_181[1:0]; // @[LZD.scala 49:47]
  assign _T_213 = _T_206[1:0]; // @[LZD.scala 49:59]
  assign _T_214 = _T_207 ? _T_212 : _T_213; // @[LZD.scala 49:35]
  assign _T_216 = {_T_209,_T_211,_T_214}; // @[Cat.scala 29:58]
  assign _T_217 = _T_155[3:0]; // @[LZD.scala 44:32]
  assign _T_218 = _T_217[3:2]; // @[LZD.scala 43:32]
  assign _T_219 = _T_218 != 2'h0; // @[LZD.scala 39:14]
  assign _T_220 = _T_218[1]; // @[LZD.scala 39:21]
  assign _T_221 = _T_218[0]; // @[LZD.scala 39:30]
  assign _T_222 = ~ _T_221; // @[LZD.scala 39:27]
  assign _T_223 = _T_220 | _T_222; // @[LZD.scala 39:25]
  assign _T_224 = {_T_219,_T_223}; // @[Cat.scala 29:58]
  assign _T_225 = _T_217[1:0]; // @[LZD.scala 44:32]
  assign _T_226 = _T_225 != 2'h0; // @[LZD.scala 39:14]
  assign _T_227 = _T_225[1]; // @[LZD.scala 39:21]
  assign _T_228 = _T_225[0]; // @[LZD.scala 39:30]
  assign _T_229 = ~ _T_228; // @[LZD.scala 39:27]
  assign _T_230 = _T_227 | _T_229; // @[LZD.scala 39:25]
  assign _T_231 = {_T_226,_T_230}; // @[Cat.scala 29:58]
  assign _T_232 = _T_224[1]; // @[Shift.scala 12:21]
  assign _T_233 = _T_231[1]; // @[Shift.scala 12:21]
  assign _T_234 = _T_232 | _T_233; // @[LZD.scala 49:16]
  assign _T_235 = ~ _T_233; // @[LZD.scala 49:27]
  assign _T_236 = _T_232 | _T_235; // @[LZD.scala 49:25]
  assign _T_237 = _T_224[0:0]; // @[LZD.scala 49:47]
  assign _T_238 = _T_231[0:0]; // @[LZD.scala 49:59]
  assign _T_239 = _T_232 ? _T_237 : _T_238; // @[LZD.scala 49:35]
  assign _T_241 = {_T_234,_T_236,_T_239}; // @[Cat.scala 29:58]
  assign _T_242 = _T_216[3]; // @[Shift.scala 12:21]
  assign _T_244 = _T_216[2:0]; // @[LZD.scala 55:32]
  assign _T_245 = _T_242 ? _T_244 : _T_241; // @[LZD.scala 55:20]
  assign _T_246 = {_T_242,_T_245}; // @[Cat.scala 29:58]
  assign _T_247 = ~ _T_246; // @[convert.scala 21:22]
  assign _T_248 = io_B[10:0]; // @[convert.scala 22:36]
  assign _T_249 = _T_247 < 4'hb; // @[Shift.scala 16:24]
  assign _T_251 = _T_247[3]; // @[Shift.scala 12:21]
  assign _T_252 = _T_248[2:0]; // @[Shift.scala 64:52]
  assign _T_254 = {_T_252,8'h0}; // @[Cat.scala 29:58]
  assign _T_255 = _T_251 ? _T_254 : _T_248; // @[Shift.scala 64:27]
  assign _T_256 = _T_247[2:0]; // @[Shift.scala 66:70]
  assign _T_257 = _T_256[2]; // @[Shift.scala 12:21]
  assign _T_258 = _T_255[6:0]; // @[Shift.scala 64:52]
  assign _T_260 = {_T_258,4'h0}; // @[Cat.scala 29:58]
  assign _T_261 = _T_257 ? _T_260 : _T_255; // @[Shift.scala 64:27]
  assign _T_262 = _T_256[1:0]; // @[Shift.scala 66:70]
  assign _T_263 = _T_262[1]; // @[Shift.scala 12:21]
  assign _T_264 = _T_261[8:0]; // @[Shift.scala 64:52]
  assign _T_266 = {_T_264,2'h0}; // @[Cat.scala 29:58]
  assign _T_267 = _T_263 ? _T_266 : _T_261; // @[Shift.scala 64:27]
  assign _T_268 = _T_262[0:0]; // @[Shift.scala 66:70]
  assign _T_270 = _T_267[9:0]; // @[Shift.scala 64:52]
  assign _T_271 = {_T_270,1'h0}; // @[Cat.scala 29:58]
  assign _T_272 = _T_268 ? _T_271 : _T_267; // @[Shift.scala 64:27]
  assign _T_273 = _T_249 ? _T_272 : 11'h0; // @[Shift.scala 16:10]
  assign _T_274 = _T_273[10:10]; // @[convert.scala 23:34]
  assign decB_fraction = _T_273[9:0]; // @[convert.scala 24:34]
  assign _T_276 = _T_152 == 1'h0; // @[convert.scala 25:26]
  assign _T_278 = _T_152 ? _T_247 : _T_246; // @[convert.scala 25:42]
  assign _T_281 = ~ _T_274; // @[convert.scala 26:67]
  assign _T_282 = _T_150 ? _T_281 : _T_274; // @[convert.scala 26:51]
  assign _T_283 = {_T_276,_T_278,_T_282}; // @[Cat.scala 29:58]
  assign _T_285 = io_B[12:0]; // @[convert.scala 29:56]
  assign _T_286 = _T_285 != 13'h0; // @[convert.scala 29:60]
  assign _T_287 = ~ _T_286; // @[convert.scala 29:41]
  assign decB_isNaR = _T_150 & _T_287; // @[convert.scala 29:39]
  assign _T_290 = _T_150 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_290 & _T_287; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_283); // @[convert.scala 32:24]
  assign aGTb = $signed(decA_scale) > $signed(decB_scale); // @[PositAdder.scala 24:32]
  assign greaterSign = aGTb ? _T_1 : _T_150; // @[PositAdder.scala 25:24]
  assign smallerSign = aGTb ? _T_150 : _T_1; // @[PositAdder.scala 26:24]
  assign greaterExp = aGTb ? $signed(decA_scale) : $signed(decB_scale); // @[PositAdder.scala 27:24]
  assign smallerExp = aGTb ? $signed(decB_scale) : $signed(decA_scale); // @[PositAdder.scala 28:24]
  assign greaterFrac = aGTb ? decA_fraction : decB_fraction; // @[PositAdder.scala 29:24]
  assign smallerFrac = aGTb ? decB_fraction : decA_fraction; // @[PositAdder.scala 30:24]
  assign smallerZero = aGTb ? decB_isZero : decA_isZero; // @[PositAdder.scala 31:24]
  assign _T_299 = $signed(greaterExp) - $signed(smallerExp); // @[PositAdder.scala 32:32]
  assign scale_diff = $signed(_T_299); // @[PositAdder.scala 32:32]
  assign _T_300 = ~ greaterSign; // @[PositAdder.scala 33:38]
  assign greaterSig = {greaterSign,_T_300,greaterFrac}; // @[Cat.scala 29:58]
  assign _T_302 = smallerSign | smallerZero; // @[PositAdder.scala 34:52]
  assign _T_303 = ~ _T_302; // @[PositAdder.scala 34:38]
  assign _T_306 = {smallerSign,_T_303,smallerFrac,3'h0}; // @[Cat.scala 29:58]
  assign _T_307 = $unsigned(scale_diff); // @[PositAdder.scala 35:68]
  assign _T_308 = _T_307 < 6'hf; // @[Shift.scala 39:24]
  assign _T_309 = _T_307[3:0]; // @[Shift.scala 40:44]
  assign _T_310 = _T_306[14:8]; // @[Shift.scala 90:30]
  assign _T_311 = _T_306[7:0]; // @[Shift.scala 90:48]
  assign _T_312 = _T_311 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_0 = {{6'd0}, _T_312}; // @[Shift.scala 90:39]
  assign _T_313 = _T_310 | _GEN_0; // @[Shift.scala 90:39]
  assign _T_314 = _T_309[3]; // @[Shift.scala 12:21]
  assign _T_315 = _T_306[14]; // @[Shift.scala 12:21]
  assign _T_317 = _T_315 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_318 = {_T_317,_T_313}; // @[Cat.scala 29:58]
  assign _T_319 = _T_314 ? _T_318 : _T_306; // @[Shift.scala 91:22]
  assign _T_320 = _T_309[2:0]; // @[Shift.scala 92:77]
  assign _T_321 = _T_319[14:4]; // @[Shift.scala 90:30]
  assign _T_322 = _T_319[3:0]; // @[Shift.scala 90:48]
  assign _T_323 = _T_322 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_1 = {{10'd0}, _T_323}; // @[Shift.scala 90:39]
  assign _T_324 = _T_321 | _GEN_1; // @[Shift.scala 90:39]
  assign _T_325 = _T_320[2]; // @[Shift.scala 12:21]
  assign _T_326 = _T_319[14]; // @[Shift.scala 12:21]
  assign _T_328 = _T_326 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_329 = {_T_328,_T_324}; // @[Cat.scala 29:58]
  assign _T_330 = _T_325 ? _T_329 : _T_319; // @[Shift.scala 91:22]
  assign _T_331 = _T_320[1:0]; // @[Shift.scala 92:77]
  assign _T_332 = _T_330[14:2]; // @[Shift.scala 90:30]
  assign _T_333 = _T_330[1:0]; // @[Shift.scala 90:48]
  assign _T_334 = _T_333 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_2 = {{12'd0}, _T_334}; // @[Shift.scala 90:39]
  assign _T_335 = _T_332 | _GEN_2; // @[Shift.scala 90:39]
  assign _T_336 = _T_331[1]; // @[Shift.scala 12:21]
  assign _T_337 = _T_330[14]; // @[Shift.scala 12:21]
  assign _T_339 = _T_337 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_340 = {_T_339,_T_335}; // @[Cat.scala 29:58]
  assign _T_341 = _T_336 ? _T_340 : _T_330; // @[Shift.scala 91:22]
  assign _T_342 = _T_331[0:0]; // @[Shift.scala 92:77]
  assign _T_343 = _T_341[14:1]; // @[Shift.scala 90:30]
  assign _T_344 = _T_341[0:0]; // @[Shift.scala 90:48]
  assign _GEN_3 = {{13'd0}, _T_344}; // @[Shift.scala 90:39]
  assign _T_346 = _T_343 | _GEN_3; // @[Shift.scala 90:39]
  assign _T_348 = _T_341[14]; // @[Shift.scala 12:21]
  assign _T_349 = {_T_348,_T_346}; // @[Cat.scala 29:58]
  assign _T_350 = _T_342 ? _T_349 : _T_341; // @[Shift.scala 91:22]
  assign _T_353 = _T_315 ? 15'h7fff : 15'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_308 ? _T_350 : _T_353; // @[Shift.scala 39:10]
  assign _T_354 = smallerSig[14:3]; // @[PositAdder.scala 36:45]
  assign rawSumSig = greaterSig + _T_354; // @[PositAdder.scala 36:32]
  assign _T_355 = _T_1 ^ _T_150; // @[PositAdder.scala 37:31]
  assign _T_356 = rawSumSig[12:12]; // @[PositAdder.scala 37:59]
  assign sumSign = _T_355 ^ _T_356; // @[PositAdder.scala 37:43]
  assign _T_357 = greaterSig + _T_354; // @[PositAdder.scala 38:48]
  assign _T_358 = smallerSig[2:0]; // @[PositAdder.scala 38:63]
  assign signSumSig = {sumSign,_T_357,_T_358}; // @[Cat.scala 29:58]
  assign _T_360 = signSumSig[15:1]; // @[PositAdder.scala 40:31]
  assign _T_361 = signSumSig[14:0]; // @[PositAdder.scala 40:66]
  assign sumXor = _T_360 ^ _T_361; // @[PositAdder.scala 40:49]
  assign _T_362 = sumXor[14:7]; // @[LZD.scala 43:32]
  assign _T_363 = _T_362[7:4]; // @[LZD.scala 43:32]
  assign _T_364 = _T_363[3:2]; // @[LZD.scala 43:32]
  assign _T_365 = _T_364 != 2'h0; // @[LZD.scala 39:14]
  assign _T_366 = _T_364[1]; // @[LZD.scala 39:21]
  assign _T_367 = _T_364[0]; // @[LZD.scala 39:30]
  assign _T_368 = ~ _T_367; // @[LZD.scala 39:27]
  assign _T_369 = _T_366 | _T_368; // @[LZD.scala 39:25]
  assign _T_370 = {_T_365,_T_369}; // @[Cat.scala 29:58]
  assign _T_371 = _T_363[1:0]; // @[LZD.scala 44:32]
  assign _T_372 = _T_371 != 2'h0; // @[LZD.scala 39:14]
  assign _T_373 = _T_371[1]; // @[LZD.scala 39:21]
  assign _T_374 = _T_371[0]; // @[LZD.scala 39:30]
  assign _T_375 = ~ _T_374; // @[LZD.scala 39:27]
  assign _T_376 = _T_373 | _T_375; // @[LZD.scala 39:25]
  assign _T_377 = {_T_372,_T_376}; // @[Cat.scala 29:58]
  assign _T_378 = _T_370[1]; // @[Shift.scala 12:21]
  assign _T_379 = _T_377[1]; // @[Shift.scala 12:21]
  assign _T_380 = _T_378 | _T_379; // @[LZD.scala 49:16]
  assign _T_381 = ~ _T_379; // @[LZD.scala 49:27]
  assign _T_382 = _T_378 | _T_381; // @[LZD.scala 49:25]
  assign _T_383 = _T_370[0:0]; // @[LZD.scala 49:47]
  assign _T_384 = _T_377[0:0]; // @[LZD.scala 49:59]
  assign _T_385 = _T_378 ? _T_383 : _T_384; // @[LZD.scala 49:35]
  assign _T_387 = {_T_380,_T_382,_T_385}; // @[Cat.scala 29:58]
  assign _T_388 = _T_362[3:0]; // @[LZD.scala 44:32]
  assign _T_389 = _T_388[3:2]; // @[LZD.scala 43:32]
  assign _T_390 = _T_389 != 2'h0; // @[LZD.scala 39:14]
  assign _T_391 = _T_389[1]; // @[LZD.scala 39:21]
  assign _T_392 = _T_389[0]; // @[LZD.scala 39:30]
  assign _T_393 = ~ _T_392; // @[LZD.scala 39:27]
  assign _T_394 = _T_391 | _T_393; // @[LZD.scala 39:25]
  assign _T_395 = {_T_390,_T_394}; // @[Cat.scala 29:58]
  assign _T_396 = _T_388[1:0]; // @[LZD.scala 44:32]
  assign _T_397 = _T_396 != 2'h0; // @[LZD.scala 39:14]
  assign _T_398 = _T_396[1]; // @[LZD.scala 39:21]
  assign _T_399 = _T_396[0]; // @[LZD.scala 39:30]
  assign _T_400 = ~ _T_399; // @[LZD.scala 39:27]
  assign _T_401 = _T_398 | _T_400; // @[LZD.scala 39:25]
  assign _T_402 = {_T_397,_T_401}; // @[Cat.scala 29:58]
  assign _T_403 = _T_395[1]; // @[Shift.scala 12:21]
  assign _T_404 = _T_402[1]; // @[Shift.scala 12:21]
  assign _T_405 = _T_403 | _T_404; // @[LZD.scala 49:16]
  assign _T_406 = ~ _T_404; // @[LZD.scala 49:27]
  assign _T_407 = _T_403 | _T_406; // @[LZD.scala 49:25]
  assign _T_408 = _T_395[0:0]; // @[LZD.scala 49:47]
  assign _T_409 = _T_402[0:0]; // @[LZD.scala 49:59]
  assign _T_410 = _T_403 ? _T_408 : _T_409; // @[LZD.scala 49:35]
  assign _T_412 = {_T_405,_T_407,_T_410}; // @[Cat.scala 29:58]
  assign _T_413 = _T_387[2]; // @[Shift.scala 12:21]
  assign _T_414 = _T_412[2]; // @[Shift.scala 12:21]
  assign _T_415 = _T_413 | _T_414; // @[LZD.scala 49:16]
  assign _T_416 = ~ _T_414; // @[LZD.scala 49:27]
  assign _T_417 = _T_413 | _T_416; // @[LZD.scala 49:25]
  assign _T_418 = _T_387[1:0]; // @[LZD.scala 49:47]
  assign _T_419 = _T_412[1:0]; // @[LZD.scala 49:59]
  assign _T_420 = _T_413 ? _T_418 : _T_419; // @[LZD.scala 49:35]
  assign _T_422 = {_T_415,_T_417,_T_420}; // @[Cat.scala 29:58]
  assign _T_423 = sumXor[6:0]; // @[LZD.scala 44:32]
  assign _T_424 = _T_423[6:3]; // @[LZD.scala 43:32]
  assign _T_425 = _T_424[3:2]; // @[LZD.scala 43:32]
  assign _T_426 = _T_425 != 2'h0; // @[LZD.scala 39:14]
  assign _T_427 = _T_425[1]; // @[LZD.scala 39:21]
  assign _T_428 = _T_425[0]; // @[LZD.scala 39:30]
  assign _T_429 = ~ _T_428; // @[LZD.scala 39:27]
  assign _T_430 = _T_427 | _T_429; // @[LZD.scala 39:25]
  assign _T_431 = {_T_426,_T_430}; // @[Cat.scala 29:58]
  assign _T_432 = _T_424[1:0]; // @[LZD.scala 44:32]
  assign _T_433 = _T_432 != 2'h0; // @[LZD.scala 39:14]
  assign _T_434 = _T_432[1]; // @[LZD.scala 39:21]
  assign _T_435 = _T_432[0]; // @[LZD.scala 39:30]
  assign _T_436 = ~ _T_435; // @[LZD.scala 39:27]
  assign _T_437 = _T_434 | _T_436; // @[LZD.scala 39:25]
  assign _T_438 = {_T_433,_T_437}; // @[Cat.scala 29:58]
  assign _T_439 = _T_431[1]; // @[Shift.scala 12:21]
  assign _T_440 = _T_438[1]; // @[Shift.scala 12:21]
  assign _T_441 = _T_439 | _T_440; // @[LZD.scala 49:16]
  assign _T_442 = ~ _T_440; // @[LZD.scala 49:27]
  assign _T_443 = _T_439 | _T_442; // @[LZD.scala 49:25]
  assign _T_444 = _T_431[0:0]; // @[LZD.scala 49:47]
  assign _T_445 = _T_438[0:0]; // @[LZD.scala 49:59]
  assign _T_446 = _T_439 ? _T_444 : _T_445; // @[LZD.scala 49:35]
  assign _T_448 = {_T_441,_T_443,_T_446}; // @[Cat.scala 29:58]
  assign _T_449 = _T_423[2:0]; // @[LZD.scala 44:32]
  assign _T_450 = _T_449[2:1]; // @[LZD.scala 43:32]
  assign _T_451 = _T_450 != 2'h0; // @[LZD.scala 39:14]
  assign _T_452 = _T_450[1]; // @[LZD.scala 39:21]
  assign _T_453 = _T_450[0]; // @[LZD.scala 39:30]
  assign _T_454 = ~ _T_453; // @[LZD.scala 39:27]
  assign _T_455 = _T_452 | _T_454; // @[LZD.scala 39:25]
  assign _T_456 = {_T_451,_T_455}; // @[Cat.scala 29:58]
  assign _T_457 = _T_449[0:0]; // @[LZD.scala 44:32]
  assign _T_459 = _T_456[1]; // @[Shift.scala 12:21]
  assign _T_461 = _T_456[0:0]; // @[LZD.scala 55:32]
  assign _T_462 = _T_459 ? _T_461 : _T_457; // @[LZD.scala 55:20]
  assign _T_463 = {_T_459,_T_462}; // @[Cat.scala 29:58]
  assign _T_464 = _T_448[2]; // @[Shift.scala 12:21]
  assign _T_466 = _T_448[1:0]; // @[LZD.scala 55:32]
  assign _T_467 = _T_464 ? _T_466 : _T_463; // @[LZD.scala 55:20]
  assign _T_468 = {_T_464,_T_467}; // @[Cat.scala 29:58]
  assign _T_469 = _T_422[3]; // @[Shift.scala 12:21]
  assign _T_471 = _T_422[2:0]; // @[LZD.scala 55:32]
  assign _T_472 = _T_469 ? _T_471 : _T_468; // @[LZD.scala 55:20]
  assign sumLZD = {_T_469,_T_472}; // @[Cat.scala 29:58]
  assign _T_473 = {1'h1,_T_469,_T_472}; // @[Cat.scala 29:58]
  assign _T_474 = $signed(_T_473); // @[PositAdder.scala 42:38]
  assign _T_476 = $signed(_T_474) + $signed(5'sh2); // @[PositAdder.scala 42:45]
  assign scaleBias = $signed(_T_476); // @[PositAdder.scala 42:45]
  assign _GEN_4 = {{1{scaleBias[4]}},scaleBias}; // @[PositAdder.scala 43:32]
  assign sumScale = $signed(greaterExp) + $signed(_GEN_4); // @[PositAdder.scala 43:32]
  assign overflow = $signed(sumScale) > $signed(7'sh18); // @[PositAdder.scala 44:30]
  assign normalShift = ~ sumLZD; // @[PositAdder.scala 45:22]
  assign _T_477 = signSumSig[13:0]; // @[PositAdder.scala 46:36]
  assign _T_478 = normalShift < 4'he; // @[Shift.scala 16:24]
  assign _T_480 = normalShift[3]; // @[Shift.scala 12:21]
  assign _T_481 = _T_477[5:0]; // @[Shift.scala 64:52]
  assign _T_483 = {_T_481,8'h0}; // @[Cat.scala 29:58]
  assign _T_484 = _T_480 ? _T_483 : _T_477; // @[Shift.scala 64:27]
  assign _T_485 = normalShift[2:0]; // @[Shift.scala 66:70]
  assign _T_486 = _T_485[2]; // @[Shift.scala 12:21]
  assign _T_487 = _T_484[9:0]; // @[Shift.scala 64:52]
  assign _T_489 = {_T_487,4'h0}; // @[Cat.scala 29:58]
  assign _T_490 = _T_486 ? _T_489 : _T_484; // @[Shift.scala 64:27]
  assign _T_491 = _T_485[1:0]; // @[Shift.scala 66:70]
  assign _T_492 = _T_491[1]; // @[Shift.scala 12:21]
  assign _T_493 = _T_490[11:0]; // @[Shift.scala 64:52]
  assign _T_495 = {_T_493,2'h0}; // @[Cat.scala 29:58]
  assign _T_496 = _T_492 ? _T_495 : _T_490; // @[Shift.scala 64:27]
  assign _T_497 = _T_491[0:0]; // @[Shift.scala 66:70]
  assign _T_499 = _T_496[12:0]; // @[Shift.scala 64:52]
  assign _T_500 = {_T_499,1'h0}; // @[Cat.scala 29:58]
  assign _T_501 = _T_497 ? _T_500 : _T_496; // @[Shift.scala 64:27]
  assign shiftSig = _T_478 ? _T_501 : 14'h0; // @[Shift.scala 16:10]
  assign _T_502 = overflow ? $signed(7'sh18) : $signed(sumScale); // @[PositAdder.scala 51:24]
  assign decS_fraction = shiftSig[13:4]; // @[PositAdder.scala 52:34]
  assign decS_isNaR = decA_isNaR | decB_isNaR; // @[PositAdder.scala 53:32]
  assign _T_505 = signSumSig != 16'h0; // @[PositAdder.scala 54:33]
  assign _T_506 = ~ _T_505; // @[PositAdder.scala 54:21]
  assign _T_507 = decA_isZero & decB_isZero; // @[PositAdder.scala 54:52]
  assign decS_isZero = _T_506 | _T_507; // @[PositAdder.scala 54:37]
  assign _T_509 = shiftSig[3:2]; // @[PositAdder.scala 55:33]
  assign _T_510 = shiftSig[1]; // @[PositAdder.scala 55:49]
  assign _T_511 = shiftSig[0]; // @[PositAdder.scala 55:63]
  assign _T_512 = _T_510 | _T_511; // @[PositAdder.scala 55:53]
  assign _GEN_5 = _T_502[5:0]; // @[PositAdder.scala 48:25 PositAdder.scala 51:18]
  assign decS_scale = $signed(_GEN_5); // @[PositAdder.scala 48:25 PositAdder.scala 51:18]
  assign _T_515 = decS_scale[0]; // @[convert.scala 46:61]
  assign _T_516 = ~ _T_515; // @[convert.scala 46:52]
  assign _T_518 = sumSign ? _T_516 : _T_515; // @[convert.scala 46:42]
  assign _T_519 = decS_scale[5:1]; // @[convert.scala 48:34]
  assign _T_520 = _T_519[4:4]; // @[convert.scala 49:36]
  assign _T_522 = ~ _T_519; // @[convert.scala 50:36]
  assign _T_523 = $signed(_T_522); // @[convert.scala 50:36]
  assign _T_524 = _T_520 ? $signed(_T_523) : $signed(_T_519); // @[convert.scala 50:28]
  assign _T_525 = _T_520 ^ sumSign; // @[convert.scala 51:31]
  assign _T_526 = ~ _T_525; // @[convert.scala 52:43]
  assign _T_530 = {_T_526,_T_525,_T_518,decS_fraction,_T_509,_T_512}; // @[Cat.scala 29:58]
  assign _T_531 = $unsigned(_T_524); // @[Shift.scala 39:17]
  assign _T_532 = _T_531 < 5'h10; // @[Shift.scala 39:24]
  assign _T_533 = _T_524[3:0]; // @[Shift.scala 40:44]
  assign _T_534 = _T_530[15:8]; // @[Shift.scala 90:30]
  assign _T_535 = _T_530[7:0]; // @[Shift.scala 90:48]
  assign _T_536 = _T_535 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_6 = {{7'd0}, _T_536}; // @[Shift.scala 90:39]
  assign _T_537 = _T_534 | _GEN_6; // @[Shift.scala 90:39]
  assign _T_538 = _T_533[3]; // @[Shift.scala 12:21]
  assign _T_539 = _T_530[15]; // @[Shift.scala 12:21]
  assign _T_541 = _T_539 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_542 = {_T_541,_T_537}; // @[Cat.scala 29:58]
  assign _T_543 = _T_538 ? _T_542 : _T_530; // @[Shift.scala 91:22]
  assign _T_544 = _T_533[2:0]; // @[Shift.scala 92:77]
  assign _T_545 = _T_543[15:4]; // @[Shift.scala 90:30]
  assign _T_546 = _T_543[3:0]; // @[Shift.scala 90:48]
  assign _T_547 = _T_546 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_7 = {{11'd0}, _T_547}; // @[Shift.scala 90:39]
  assign _T_548 = _T_545 | _GEN_7; // @[Shift.scala 90:39]
  assign _T_549 = _T_544[2]; // @[Shift.scala 12:21]
  assign _T_550 = _T_543[15]; // @[Shift.scala 12:21]
  assign _T_552 = _T_550 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_553 = {_T_552,_T_548}; // @[Cat.scala 29:58]
  assign _T_554 = _T_549 ? _T_553 : _T_543; // @[Shift.scala 91:22]
  assign _T_555 = _T_544[1:0]; // @[Shift.scala 92:77]
  assign _T_556 = _T_554[15:2]; // @[Shift.scala 90:30]
  assign _T_557 = _T_554[1:0]; // @[Shift.scala 90:48]
  assign _T_558 = _T_557 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_8 = {{13'd0}, _T_558}; // @[Shift.scala 90:39]
  assign _T_559 = _T_556 | _GEN_8; // @[Shift.scala 90:39]
  assign _T_560 = _T_555[1]; // @[Shift.scala 12:21]
  assign _T_561 = _T_554[15]; // @[Shift.scala 12:21]
  assign _T_563 = _T_561 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_564 = {_T_563,_T_559}; // @[Cat.scala 29:58]
  assign _T_565 = _T_560 ? _T_564 : _T_554; // @[Shift.scala 91:22]
  assign _T_566 = _T_555[0:0]; // @[Shift.scala 92:77]
  assign _T_567 = _T_565[15:1]; // @[Shift.scala 90:30]
  assign _T_568 = _T_565[0:0]; // @[Shift.scala 90:48]
  assign _GEN_9 = {{14'd0}, _T_568}; // @[Shift.scala 90:39]
  assign _T_570 = _T_567 | _GEN_9; // @[Shift.scala 90:39]
  assign _T_572 = _T_565[15]; // @[Shift.scala 12:21]
  assign _T_573 = {_T_572,_T_570}; // @[Cat.scala 29:58]
  assign _T_574 = _T_566 ? _T_573 : _T_565; // @[Shift.scala 91:22]
  assign _T_577 = _T_539 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_578 = _T_532 ? _T_574 : _T_577; // @[Shift.scala 39:10]
  assign _T_579 = _T_578[3]; // @[convert.scala 55:31]
  assign _T_580 = _T_578[2]; // @[convert.scala 56:31]
  assign _T_581 = _T_578[1]; // @[convert.scala 57:31]
  assign _T_582 = _T_578[0]; // @[convert.scala 58:31]
  assign _T_583 = _T_578[15:3]; // @[convert.scala 59:69]
  assign _T_584 = _T_583 != 13'h0; // @[convert.scala 59:81]
  assign _T_585 = ~ _T_584; // @[convert.scala 59:50]
  assign _T_587 = _T_583 == 13'h1fff; // @[convert.scala 60:81]
  assign _T_588 = _T_579 | _T_581; // @[convert.scala 61:44]
  assign _T_589 = _T_588 | _T_582; // @[convert.scala 61:52]
  assign _T_590 = _T_580 & _T_589; // @[convert.scala 61:36]
  assign _T_591 = ~ _T_587; // @[convert.scala 62:63]
  assign _T_592 = _T_591 & _T_590; // @[convert.scala 62:103]
  assign _T_593 = _T_585 | _T_592; // @[convert.scala 62:60]
  assign _GEN_10 = {{12'd0}, _T_593}; // @[convert.scala 63:56]
  assign _T_596 = _T_583 + _GEN_10; // @[convert.scala 63:56]
  assign _T_597 = {sumSign,_T_596}; // @[Cat.scala 29:58]
  assign _T_599 = decS_isZero ? 14'h0 : _T_597; // @[Mux.scala 87:16]
  assign io_S = decS_isNaR ? 14'h2000 : _T_599; // @[PositAdder.scala 57:8]
endmodule
