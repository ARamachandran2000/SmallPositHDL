module PositFMA16_1(
  input         clock,
  input         reset,
  input         io_inValid,
  input  [1:0]  io_fmaOp,
  input  [15:0] io_A,
  input  [15:0] io_B,
  input  [15:0] io_C,
  output [15:0] io_F,
  output        io_outValid
);
  wire  _T; // @[PositFMA.scala 47:36]
  wire [15:0] _T_2; // @[Bitwise.scala 71:12]
  wire [15:0] _T_3; // @[PositFMA.scala 47:41]
  wire [15:0] _GEN_10; // @[PositFMA.scala 47:49]
  wire [15:0] realA; // @[PositFMA.scala 47:49]
  wire  _T_6; // @[PositFMA.scala 48:36]
  wire [15:0] _T_8; // @[Bitwise.scala 71:12]
  wire [15:0] _T_9; // @[PositFMA.scala 48:41]
  wire [15:0] _GEN_11; // @[PositFMA.scala 48:49]
  wire [15:0] realC; // @[PositFMA.scala 48:49]
  wire  _T_13; // @[convert.scala 18:24]
  wire  _T_14; // @[convert.scala 18:40]
  wire  _T_15; // @[convert.scala 18:36]
  wire [13:0] _T_16; // @[convert.scala 19:24]
  wire [13:0] _T_17; // @[convert.scala 19:43]
  wire [13:0] _T_18; // @[convert.scala 19:39]
  wire [7:0] _T_19; // @[LZD.scala 43:32]
  wire [3:0] _T_20; // @[LZD.scala 43:32]
  wire [1:0] _T_21; // @[LZD.scala 43:32]
  wire  _T_22; // @[LZD.scala 39:14]
  wire  _T_23; // @[LZD.scala 39:21]
  wire  _T_24; // @[LZD.scala 39:30]
  wire  _T_25; // @[LZD.scala 39:27]
  wire  _T_26; // @[LZD.scala 39:25]
  wire [1:0] _T_27; // @[Cat.scala 29:58]
  wire [1:0] _T_28; // @[LZD.scala 44:32]
  wire  _T_29; // @[LZD.scala 39:14]
  wire  _T_30; // @[LZD.scala 39:21]
  wire  _T_31; // @[LZD.scala 39:30]
  wire  _T_32; // @[LZD.scala 39:27]
  wire  _T_33; // @[LZD.scala 39:25]
  wire [1:0] _T_34; // @[Cat.scala 29:58]
  wire  _T_35; // @[Shift.scala 12:21]
  wire  _T_36; // @[Shift.scala 12:21]
  wire  _T_37; // @[LZD.scala 49:16]
  wire  _T_38; // @[LZD.scala 49:27]
  wire  _T_39; // @[LZD.scala 49:25]
  wire  _T_40; // @[LZD.scala 49:47]
  wire  _T_41; // @[LZD.scala 49:59]
  wire  _T_42; // @[LZD.scala 49:35]
  wire [2:0] _T_44; // @[Cat.scala 29:58]
  wire [3:0] _T_45; // @[LZD.scala 44:32]
  wire [1:0] _T_46; // @[LZD.scala 43:32]
  wire  _T_47; // @[LZD.scala 39:14]
  wire  _T_48; // @[LZD.scala 39:21]
  wire  _T_49; // @[LZD.scala 39:30]
  wire  _T_50; // @[LZD.scala 39:27]
  wire  _T_51; // @[LZD.scala 39:25]
  wire [1:0] _T_52; // @[Cat.scala 29:58]
  wire [1:0] _T_53; // @[LZD.scala 44:32]
  wire  _T_54; // @[LZD.scala 39:14]
  wire  _T_55; // @[LZD.scala 39:21]
  wire  _T_56; // @[LZD.scala 39:30]
  wire  _T_57; // @[LZD.scala 39:27]
  wire  _T_58; // @[LZD.scala 39:25]
  wire [1:0] _T_59; // @[Cat.scala 29:58]
  wire  _T_60; // @[Shift.scala 12:21]
  wire  _T_61; // @[Shift.scala 12:21]
  wire  _T_62; // @[LZD.scala 49:16]
  wire  _T_63; // @[LZD.scala 49:27]
  wire  _T_64; // @[LZD.scala 49:25]
  wire  _T_65; // @[LZD.scala 49:47]
  wire  _T_66; // @[LZD.scala 49:59]
  wire  _T_67; // @[LZD.scala 49:35]
  wire [2:0] _T_69; // @[Cat.scala 29:58]
  wire  _T_70; // @[Shift.scala 12:21]
  wire  _T_71; // @[Shift.scala 12:21]
  wire  _T_72; // @[LZD.scala 49:16]
  wire  _T_73; // @[LZD.scala 49:27]
  wire  _T_74; // @[LZD.scala 49:25]
  wire [1:0] _T_75; // @[LZD.scala 49:47]
  wire [1:0] _T_76; // @[LZD.scala 49:59]
  wire [1:0] _T_77; // @[LZD.scala 49:35]
  wire [3:0] _T_79; // @[Cat.scala 29:58]
  wire [5:0] _T_80; // @[LZD.scala 44:32]
  wire [3:0] _T_81; // @[LZD.scala 43:32]
  wire [1:0] _T_82; // @[LZD.scala 43:32]
  wire  _T_83; // @[LZD.scala 39:14]
  wire  _T_84; // @[LZD.scala 39:21]
  wire  _T_85; // @[LZD.scala 39:30]
  wire  _T_86; // @[LZD.scala 39:27]
  wire  _T_87; // @[LZD.scala 39:25]
  wire [1:0] _T_88; // @[Cat.scala 29:58]
  wire [1:0] _T_89; // @[LZD.scala 44:32]
  wire  _T_90; // @[LZD.scala 39:14]
  wire  _T_91; // @[LZD.scala 39:21]
  wire  _T_92; // @[LZD.scala 39:30]
  wire  _T_93; // @[LZD.scala 39:27]
  wire  _T_94; // @[LZD.scala 39:25]
  wire [1:0] _T_95; // @[Cat.scala 29:58]
  wire  _T_96; // @[Shift.scala 12:21]
  wire  _T_97; // @[Shift.scala 12:21]
  wire  _T_98; // @[LZD.scala 49:16]
  wire  _T_99; // @[LZD.scala 49:27]
  wire  _T_100; // @[LZD.scala 49:25]
  wire  _T_101; // @[LZD.scala 49:47]
  wire  _T_102; // @[LZD.scala 49:59]
  wire  _T_103; // @[LZD.scala 49:35]
  wire [2:0] _T_105; // @[Cat.scala 29:58]
  wire [1:0] _T_106; // @[LZD.scala 44:32]
  wire  _T_107; // @[LZD.scala 39:14]
  wire  _T_108; // @[LZD.scala 39:21]
  wire  _T_109; // @[LZD.scala 39:30]
  wire  _T_110; // @[LZD.scala 39:27]
  wire  _T_111; // @[LZD.scala 39:25]
  wire [1:0] _T_112; // @[Cat.scala 29:58]
  wire  _T_113; // @[Shift.scala 12:21]
  wire [1:0] _T_115; // @[LZD.scala 55:32]
  wire [1:0] _T_116; // @[LZD.scala 55:20]
  wire [2:0] _T_117; // @[Cat.scala 29:58]
  wire  _T_118; // @[Shift.scala 12:21]
  wire [2:0] _T_120; // @[LZD.scala 55:32]
  wire [2:0] _T_121; // @[LZD.scala 55:20]
  wire [3:0] _T_122; // @[Cat.scala 29:58]
  wire [3:0] _T_123; // @[convert.scala 21:22]
  wire [12:0] _T_124; // @[convert.scala 22:36]
  wire  _T_125; // @[Shift.scala 16:24]
  wire  _T_127; // @[Shift.scala 12:21]
  wire [4:0] _T_128; // @[Shift.scala 64:52]
  wire [12:0] _T_130; // @[Cat.scala 29:58]
  wire [12:0] _T_131; // @[Shift.scala 64:27]
  wire [2:0] _T_132; // @[Shift.scala 66:70]
  wire  _T_133; // @[Shift.scala 12:21]
  wire [8:0] _T_134; // @[Shift.scala 64:52]
  wire [12:0] _T_136; // @[Cat.scala 29:58]
  wire [12:0] _T_137; // @[Shift.scala 64:27]
  wire [1:0] _T_138; // @[Shift.scala 66:70]
  wire  _T_139; // @[Shift.scala 12:21]
  wire [10:0] _T_140; // @[Shift.scala 64:52]
  wire [12:0] _T_142; // @[Cat.scala 29:58]
  wire [12:0] _T_143; // @[Shift.scala 64:27]
  wire  _T_144; // @[Shift.scala 66:70]
  wire [11:0] _T_146; // @[Shift.scala 64:52]
  wire [12:0] _T_147; // @[Cat.scala 29:58]
  wire [12:0] _T_148; // @[Shift.scala 64:27]
  wire [12:0] _T_149; // @[Shift.scala 16:10]
  wire  _T_150; // @[convert.scala 23:34]
  wire [11:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_152; // @[convert.scala 25:26]
  wire [3:0] _T_154; // @[convert.scala 25:42]
  wire  _T_157; // @[convert.scala 26:67]
  wire  _T_158; // @[convert.scala 26:51]
  wire [5:0] _T_159; // @[Cat.scala 29:58]
  wire [14:0] _T_161; // @[convert.scala 29:56]
  wire  _T_162; // @[convert.scala 29:60]
  wire  _T_163; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_166; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [5:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_175; // @[convert.scala 18:24]
  wire  _T_176; // @[convert.scala 18:40]
  wire  _T_177; // @[convert.scala 18:36]
  wire [13:0] _T_178; // @[convert.scala 19:24]
  wire [13:0] _T_179; // @[convert.scala 19:43]
  wire [13:0] _T_180; // @[convert.scala 19:39]
  wire [7:0] _T_181; // @[LZD.scala 43:32]
  wire [3:0] _T_182; // @[LZD.scala 43:32]
  wire [1:0] _T_183; // @[LZD.scala 43:32]
  wire  _T_184; // @[LZD.scala 39:14]
  wire  _T_185; // @[LZD.scala 39:21]
  wire  _T_186; // @[LZD.scala 39:30]
  wire  _T_187; // @[LZD.scala 39:27]
  wire  _T_188; // @[LZD.scala 39:25]
  wire [1:0] _T_189; // @[Cat.scala 29:58]
  wire [1:0] _T_190; // @[LZD.scala 44:32]
  wire  _T_191; // @[LZD.scala 39:14]
  wire  _T_192; // @[LZD.scala 39:21]
  wire  _T_193; // @[LZD.scala 39:30]
  wire  _T_194; // @[LZD.scala 39:27]
  wire  _T_195; // @[LZD.scala 39:25]
  wire [1:0] _T_196; // @[Cat.scala 29:58]
  wire  _T_197; // @[Shift.scala 12:21]
  wire  _T_198; // @[Shift.scala 12:21]
  wire  _T_199; // @[LZD.scala 49:16]
  wire  _T_200; // @[LZD.scala 49:27]
  wire  _T_201; // @[LZD.scala 49:25]
  wire  _T_202; // @[LZD.scala 49:47]
  wire  _T_203; // @[LZD.scala 49:59]
  wire  _T_204; // @[LZD.scala 49:35]
  wire [2:0] _T_206; // @[Cat.scala 29:58]
  wire [3:0] _T_207; // @[LZD.scala 44:32]
  wire [1:0] _T_208; // @[LZD.scala 43:32]
  wire  _T_209; // @[LZD.scala 39:14]
  wire  _T_210; // @[LZD.scala 39:21]
  wire  _T_211; // @[LZD.scala 39:30]
  wire  _T_212; // @[LZD.scala 39:27]
  wire  _T_213; // @[LZD.scala 39:25]
  wire [1:0] _T_214; // @[Cat.scala 29:58]
  wire [1:0] _T_215; // @[LZD.scala 44:32]
  wire  _T_216; // @[LZD.scala 39:14]
  wire  _T_217; // @[LZD.scala 39:21]
  wire  _T_218; // @[LZD.scala 39:30]
  wire  _T_219; // @[LZD.scala 39:27]
  wire  _T_220; // @[LZD.scala 39:25]
  wire [1:0] _T_221; // @[Cat.scala 29:58]
  wire  _T_222; // @[Shift.scala 12:21]
  wire  _T_223; // @[Shift.scala 12:21]
  wire  _T_224; // @[LZD.scala 49:16]
  wire  _T_225; // @[LZD.scala 49:27]
  wire  _T_226; // @[LZD.scala 49:25]
  wire  _T_227; // @[LZD.scala 49:47]
  wire  _T_228; // @[LZD.scala 49:59]
  wire  _T_229; // @[LZD.scala 49:35]
  wire [2:0] _T_231; // @[Cat.scala 29:58]
  wire  _T_232; // @[Shift.scala 12:21]
  wire  _T_233; // @[Shift.scala 12:21]
  wire  _T_234; // @[LZD.scala 49:16]
  wire  _T_235; // @[LZD.scala 49:27]
  wire  _T_236; // @[LZD.scala 49:25]
  wire [1:0] _T_237; // @[LZD.scala 49:47]
  wire [1:0] _T_238; // @[LZD.scala 49:59]
  wire [1:0] _T_239; // @[LZD.scala 49:35]
  wire [3:0] _T_241; // @[Cat.scala 29:58]
  wire [5:0] _T_242; // @[LZD.scala 44:32]
  wire [3:0] _T_243; // @[LZD.scala 43:32]
  wire [1:0] _T_244; // @[LZD.scala 43:32]
  wire  _T_245; // @[LZD.scala 39:14]
  wire  _T_246; // @[LZD.scala 39:21]
  wire  _T_247; // @[LZD.scala 39:30]
  wire  _T_248; // @[LZD.scala 39:27]
  wire  _T_249; // @[LZD.scala 39:25]
  wire [1:0] _T_250; // @[Cat.scala 29:58]
  wire [1:0] _T_251; // @[LZD.scala 44:32]
  wire  _T_252; // @[LZD.scala 39:14]
  wire  _T_253; // @[LZD.scala 39:21]
  wire  _T_254; // @[LZD.scala 39:30]
  wire  _T_255; // @[LZD.scala 39:27]
  wire  _T_256; // @[LZD.scala 39:25]
  wire [1:0] _T_257; // @[Cat.scala 29:58]
  wire  _T_258; // @[Shift.scala 12:21]
  wire  _T_259; // @[Shift.scala 12:21]
  wire  _T_260; // @[LZD.scala 49:16]
  wire  _T_261; // @[LZD.scala 49:27]
  wire  _T_262; // @[LZD.scala 49:25]
  wire  _T_263; // @[LZD.scala 49:47]
  wire  _T_264; // @[LZD.scala 49:59]
  wire  _T_265; // @[LZD.scala 49:35]
  wire [2:0] _T_267; // @[Cat.scala 29:58]
  wire [1:0] _T_268; // @[LZD.scala 44:32]
  wire  _T_269; // @[LZD.scala 39:14]
  wire  _T_270; // @[LZD.scala 39:21]
  wire  _T_271; // @[LZD.scala 39:30]
  wire  _T_272; // @[LZD.scala 39:27]
  wire  _T_273; // @[LZD.scala 39:25]
  wire [1:0] _T_274; // @[Cat.scala 29:58]
  wire  _T_275; // @[Shift.scala 12:21]
  wire [1:0] _T_277; // @[LZD.scala 55:32]
  wire [1:0] _T_278; // @[LZD.scala 55:20]
  wire [2:0] _T_279; // @[Cat.scala 29:58]
  wire  _T_280; // @[Shift.scala 12:21]
  wire [2:0] _T_282; // @[LZD.scala 55:32]
  wire [2:0] _T_283; // @[LZD.scala 55:20]
  wire [3:0] _T_284; // @[Cat.scala 29:58]
  wire [3:0] _T_285; // @[convert.scala 21:22]
  wire [12:0] _T_286; // @[convert.scala 22:36]
  wire  _T_287; // @[Shift.scala 16:24]
  wire  _T_289; // @[Shift.scala 12:21]
  wire [4:0] _T_290; // @[Shift.scala 64:52]
  wire [12:0] _T_292; // @[Cat.scala 29:58]
  wire [12:0] _T_293; // @[Shift.scala 64:27]
  wire [2:0] _T_294; // @[Shift.scala 66:70]
  wire  _T_295; // @[Shift.scala 12:21]
  wire [8:0] _T_296; // @[Shift.scala 64:52]
  wire [12:0] _T_298; // @[Cat.scala 29:58]
  wire [12:0] _T_299; // @[Shift.scala 64:27]
  wire [1:0] _T_300; // @[Shift.scala 66:70]
  wire  _T_301; // @[Shift.scala 12:21]
  wire [10:0] _T_302; // @[Shift.scala 64:52]
  wire [12:0] _T_304; // @[Cat.scala 29:58]
  wire [12:0] _T_305; // @[Shift.scala 64:27]
  wire  _T_306; // @[Shift.scala 66:70]
  wire [11:0] _T_308; // @[Shift.scala 64:52]
  wire [12:0] _T_309; // @[Cat.scala 29:58]
  wire [12:0] _T_310; // @[Shift.scala 64:27]
  wire [12:0] _T_311; // @[Shift.scala 16:10]
  wire  _T_312; // @[convert.scala 23:34]
  wire [11:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_314; // @[convert.scala 25:26]
  wire [3:0] _T_316; // @[convert.scala 25:42]
  wire  _T_319; // @[convert.scala 26:67]
  wire  _T_320; // @[convert.scala 26:51]
  wire [5:0] _T_321; // @[Cat.scala 29:58]
  wire [14:0] _T_323; // @[convert.scala 29:56]
  wire  _T_324; // @[convert.scala 29:60]
  wire  _T_325; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_328; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [5:0] decB_scale; // @[convert.scala 32:24]
  wire  _T_337; // @[convert.scala 18:24]
  wire  _T_338; // @[convert.scala 18:40]
  wire  _T_339; // @[convert.scala 18:36]
  wire [13:0] _T_340; // @[convert.scala 19:24]
  wire [13:0] _T_341; // @[convert.scala 19:43]
  wire [13:0] _T_342; // @[convert.scala 19:39]
  wire [7:0] _T_343; // @[LZD.scala 43:32]
  wire [3:0] _T_344; // @[LZD.scala 43:32]
  wire [1:0] _T_345; // @[LZD.scala 43:32]
  wire  _T_346; // @[LZD.scala 39:14]
  wire  _T_347; // @[LZD.scala 39:21]
  wire  _T_348; // @[LZD.scala 39:30]
  wire  _T_349; // @[LZD.scala 39:27]
  wire  _T_350; // @[LZD.scala 39:25]
  wire [1:0] _T_351; // @[Cat.scala 29:58]
  wire [1:0] _T_352; // @[LZD.scala 44:32]
  wire  _T_353; // @[LZD.scala 39:14]
  wire  _T_354; // @[LZD.scala 39:21]
  wire  _T_355; // @[LZD.scala 39:30]
  wire  _T_356; // @[LZD.scala 39:27]
  wire  _T_357; // @[LZD.scala 39:25]
  wire [1:0] _T_358; // @[Cat.scala 29:58]
  wire  _T_359; // @[Shift.scala 12:21]
  wire  _T_360; // @[Shift.scala 12:21]
  wire  _T_361; // @[LZD.scala 49:16]
  wire  _T_362; // @[LZD.scala 49:27]
  wire  _T_363; // @[LZD.scala 49:25]
  wire  _T_364; // @[LZD.scala 49:47]
  wire  _T_365; // @[LZD.scala 49:59]
  wire  _T_366; // @[LZD.scala 49:35]
  wire [2:0] _T_368; // @[Cat.scala 29:58]
  wire [3:0] _T_369; // @[LZD.scala 44:32]
  wire [1:0] _T_370; // @[LZD.scala 43:32]
  wire  _T_371; // @[LZD.scala 39:14]
  wire  _T_372; // @[LZD.scala 39:21]
  wire  _T_373; // @[LZD.scala 39:30]
  wire  _T_374; // @[LZD.scala 39:27]
  wire  _T_375; // @[LZD.scala 39:25]
  wire [1:0] _T_376; // @[Cat.scala 29:58]
  wire [1:0] _T_377; // @[LZD.scala 44:32]
  wire  _T_378; // @[LZD.scala 39:14]
  wire  _T_379; // @[LZD.scala 39:21]
  wire  _T_380; // @[LZD.scala 39:30]
  wire  _T_381; // @[LZD.scala 39:27]
  wire  _T_382; // @[LZD.scala 39:25]
  wire [1:0] _T_383; // @[Cat.scala 29:58]
  wire  _T_384; // @[Shift.scala 12:21]
  wire  _T_385; // @[Shift.scala 12:21]
  wire  _T_386; // @[LZD.scala 49:16]
  wire  _T_387; // @[LZD.scala 49:27]
  wire  _T_388; // @[LZD.scala 49:25]
  wire  _T_389; // @[LZD.scala 49:47]
  wire  _T_390; // @[LZD.scala 49:59]
  wire  _T_391; // @[LZD.scala 49:35]
  wire [2:0] _T_393; // @[Cat.scala 29:58]
  wire  _T_394; // @[Shift.scala 12:21]
  wire  _T_395; // @[Shift.scala 12:21]
  wire  _T_396; // @[LZD.scala 49:16]
  wire  _T_397; // @[LZD.scala 49:27]
  wire  _T_398; // @[LZD.scala 49:25]
  wire [1:0] _T_399; // @[LZD.scala 49:47]
  wire [1:0] _T_400; // @[LZD.scala 49:59]
  wire [1:0] _T_401; // @[LZD.scala 49:35]
  wire [3:0] _T_403; // @[Cat.scala 29:58]
  wire [5:0] _T_404; // @[LZD.scala 44:32]
  wire [3:0] _T_405; // @[LZD.scala 43:32]
  wire [1:0] _T_406; // @[LZD.scala 43:32]
  wire  _T_407; // @[LZD.scala 39:14]
  wire  _T_408; // @[LZD.scala 39:21]
  wire  _T_409; // @[LZD.scala 39:30]
  wire  _T_410; // @[LZD.scala 39:27]
  wire  _T_411; // @[LZD.scala 39:25]
  wire [1:0] _T_412; // @[Cat.scala 29:58]
  wire [1:0] _T_413; // @[LZD.scala 44:32]
  wire  _T_414; // @[LZD.scala 39:14]
  wire  _T_415; // @[LZD.scala 39:21]
  wire  _T_416; // @[LZD.scala 39:30]
  wire  _T_417; // @[LZD.scala 39:27]
  wire  _T_418; // @[LZD.scala 39:25]
  wire [1:0] _T_419; // @[Cat.scala 29:58]
  wire  _T_420; // @[Shift.scala 12:21]
  wire  _T_421; // @[Shift.scala 12:21]
  wire  _T_422; // @[LZD.scala 49:16]
  wire  _T_423; // @[LZD.scala 49:27]
  wire  _T_424; // @[LZD.scala 49:25]
  wire  _T_425; // @[LZD.scala 49:47]
  wire  _T_426; // @[LZD.scala 49:59]
  wire  _T_427; // @[LZD.scala 49:35]
  wire [2:0] _T_429; // @[Cat.scala 29:58]
  wire [1:0] _T_430; // @[LZD.scala 44:32]
  wire  _T_431; // @[LZD.scala 39:14]
  wire  _T_432; // @[LZD.scala 39:21]
  wire  _T_433; // @[LZD.scala 39:30]
  wire  _T_434; // @[LZD.scala 39:27]
  wire  _T_435; // @[LZD.scala 39:25]
  wire [1:0] _T_436; // @[Cat.scala 29:58]
  wire  _T_437; // @[Shift.scala 12:21]
  wire [1:0] _T_439; // @[LZD.scala 55:32]
  wire [1:0] _T_440; // @[LZD.scala 55:20]
  wire [2:0] _T_441; // @[Cat.scala 29:58]
  wire  _T_442; // @[Shift.scala 12:21]
  wire [2:0] _T_444; // @[LZD.scala 55:32]
  wire [2:0] _T_445; // @[LZD.scala 55:20]
  wire [3:0] _T_446; // @[Cat.scala 29:58]
  wire [3:0] _T_447; // @[convert.scala 21:22]
  wire [12:0] _T_448; // @[convert.scala 22:36]
  wire  _T_449; // @[Shift.scala 16:24]
  wire  _T_451; // @[Shift.scala 12:21]
  wire [4:0] _T_452; // @[Shift.scala 64:52]
  wire [12:0] _T_454; // @[Cat.scala 29:58]
  wire [12:0] _T_455; // @[Shift.scala 64:27]
  wire [2:0] _T_456; // @[Shift.scala 66:70]
  wire  _T_457; // @[Shift.scala 12:21]
  wire [8:0] _T_458; // @[Shift.scala 64:52]
  wire [12:0] _T_460; // @[Cat.scala 29:58]
  wire [12:0] _T_461; // @[Shift.scala 64:27]
  wire [1:0] _T_462; // @[Shift.scala 66:70]
  wire  _T_463; // @[Shift.scala 12:21]
  wire [10:0] _T_464; // @[Shift.scala 64:52]
  wire [12:0] _T_466; // @[Cat.scala 29:58]
  wire [12:0] _T_467; // @[Shift.scala 64:27]
  wire  _T_468; // @[Shift.scala 66:70]
  wire [11:0] _T_470; // @[Shift.scala 64:52]
  wire [12:0] _T_471; // @[Cat.scala 29:58]
  wire [12:0] _T_472; // @[Shift.scala 64:27]
  wire [12:0] _T_473; // @[Shift.scala 16:10]
  wire  _T_474; // @[convert.scala 23:34]
  wire [11:0] decC_fraction; // @[convert.scala 24:34]
  wire  _T_476; // @[convert.scala 25:26]
  wire [3:0] _T_478; // @[convert.scala 25:42]
  wire  _T_481; // @[convert.scala 26:67]
  wire  _T_482; // @[convert.scala 26:51]
  wire [5:0] _T_483; // @[Cat.scala 29:58]
  wire [14:0] _T_485; // @[convert.scala 29:56]
  wire  _T_486; // @[convert.scala 29:60]
  wire  _T_487; // @[convert.scala 29:41]
  wire  decC_isNaR; // @[convert.scala 29:39]
  wire  _T_490; // @[convert.scala 30:19]
  wire  decC_isZero; // @[convert.scala 30:41]
  wire [5:0] decC_scale; // @[convert.scala 32:24]
  wire  _T_498; // @[PositFMA.scala 58:30]
  wire  outIsNaR; // @[PositFMA.scala 58:44]
  wire  _T_499; // @[PositFMA.scala 59:34]
  wire  _T_500; // @[PositFMA.scala 59:47]
  wire  _T_501; // @[PositFMA.scala 59:45]
  wire [13:0] _T_503; // @[Cat.scala 29:58]
  wire [13:0] sigA; // @[PositFMA.scala 59:76]
  wire  _T_504; // @[PositFMA.scala 60:34]
  wire  _T_505; // @[PositFMA.scala 60:47]
  wire  _T_506; // @[PositFMA.scala 60:45]
  wire [13:0] _T_508; // @[Cat.scala 29:58]
  wire [13:0] sigB; // @[PositFMA.scala 60:76]
  wire [27:0] _T_509; // @[PositFMA.scala 61:25]
  wire [27:0] sigP; // @[PositFMA.scala 61:33]
  wire [1:0] head2; // @[PositFMA.scala 62:28]
  wire  _T_510; // @[PositFMA.scala 63:31]
  wire  _T_511; // @[PositFMA.scala 63:25]
  wire  _T_512; // @[PositFMA.scala 63:42]
  wire  addTwo; // @[PositFMA.scala 63:35]
  wire  _T_513; // @[PositFMA.scala 65:23]
  wire  _T_514; // @[PositFMA.scala 65:49]
  wire  addOne; // @[PositFMA.scala 65:43]
  wire [1:0] _T_515; // @[Cat.scala 29:58]
  wire [2:0] expBias; // @[PositFMA.scala 66:39]
  wire  mulSign; // @[PositFMA.scala 67:28]
  wire [6:0] _T_516; // @[PositFMA.scala 69:30]
  wire [6:0] _GEN_12; // @[PositFMA.scala 69:44]
  wire [6:0] _T_518; // @[PositFMA.scala 69:44]
  wire [6:0] mulScale; // @[PositFMA.scala 69:44]
  wire [25:0] _T_519; // @[PositFMA.scala 72:29]
  wire [24:0] _T_520; // @[PositFMA.scala 73:29]
  wire [25:0] _T_521; // @[PositFMA.scala 73:48]
  wire [25:0] mulSigTmp; // @[PositFMA.scala 70:22]
  wire  _T_523; // @[PositFMA.scala 77:39]
  wire  _T_524; // @[PositFMA.scala 77:43]
  wire [24:0] _T_525; // @[PositFMA.scala 78:39]
  wire [26:0] mulSig; // @[Cat.scala 29:58]
  reg  outIsNaR_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg [26:0] mulSig_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg [11:0] addFrac_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [6:0] mulScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [5:0] addScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  addSign_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  addZero_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  inValid_phase2; // @[Valid.scala 117:22]
  reg [31:0] _RAND_7;
  wire  _T_551; // @[PositFMA.scala 107:29]
  wire  _T_552; // @[PositFMA.scala 107:47]
  wire  _T_553; // @[PositFMA.scala 107:45]
  wire [26:0] extAddSig; // @[Cat.scala 29:58]
  wire [6:0] _GEN_13; // @[PositFMA.scala 111:39]
  wire  mulGreater; // @[PositFMA.scala 111:39]
  wire [6:0] greaterScale; // @[PositFMA.scala 112:26]
  wire [6:0] smallerScale; // @[PositFMA.scala 113:26]
  wire [6:0] _T_557; // @[PositFMA.scala 114:36]
  wire [6:0] scaleDiff; // @[PositFMA.scala 114:36]
  wire [26:0] greaterSig; // @[PositFMA.scala 115:26]
  wire [26:0] smallerSigTmp; // @[PositFMA.scala 116:26]
  wire [6:0] _T_558; // @[PositFMA.scala 117:69]
  wire  _T_559; // @[Shift.scala 39:24]
  wire [4:0] _T_560; // @[Shift.scala 40:44]
  wire [10:0] _T_561; // @[Shift.scala 90:30]
  wire [15:0] _T_562; // @[Shift.scala 90:48]
  wire  _T_563; // @[Shift.scala 90:57]
  wire [10:0] _GEN_14; // @[Shift.scala 90:39]
  wire [10:0] _T_564; // @[Shift.scala 90:39]
  wire  _T_565; // @[Shift.scala 12:21]
  wire  _T_566; // @[Shift.scala 12:21]
  wire [15:0] _T_568; // @[Bitwise.scala 71:12]
  wire [26:0] _T_569; // @[Cat.scala 29:58]
  wire [26:0] _T_570; // @[Shift.scala 91:22]
  wire [3:0] _T_571; // @[Shift.scala 92:77]
  wire [18:0] _T_572; // @[Shift.scala 90:30]
  wire [7:0] _T_573; // @[Shift.scala 90:48]
  wire  _T_574; // @[Shift.scala 90:57]
  wire [18:0] _GEN_15; // @[Shift.scala 90:39]
  wire [18:0] _T_575; // @[Shift.scala 90:39]
  wire  _T_576; // @[Shift.scala 12:21]
  wire  _T_577; // @[Shift.scala 12:21]
  wire [7:0] _T_579; // @[Bitwise.scala 71:12]
  wire [26:0] _T_580; // @[Cat.scala 29:58]
  wire [26:0] _T_581; // @[Shift.scala 91:22]
  wire [2:0] _T_582; // @[Shift.scala 92:77]
  wire [22:0] _T_583; // @[Shift.scala 90:30]
  wire [3:0] _T_584; // @[Shift.scala 90:48]
  wire  _T_585; // @[Shift.scala 90:57]
  wire [22:0] _GEN_16; // @[Shift.scala 90:39]
  wire [22:0] _T_586; // @[Shift.scala 90:39]
  wire  _T_587; // @[Shift.scala 12:21]
  wire  _T_588; // @[Shift.scala 12:21]
  wire [3:0] _T_590; // @[Bitwise.scala 71:12]
  wire [26:0] _T_591; // @[Cat.scala 29:58]
  wire [26:0] _T_592; // @[Shift.scala 91:22]
  wire [1:0] _T_593; // @[Shift.scala 92:77]
  wire [24:0] _T_594; // @[Shift.scala 90:30]
  wire [1:0] _T_595; // @[Shift.scala 90:48]
  wire  _T_596; // @[Shift.scala 90:57]
  wire [24:0] _GEN_17; // @[Shift.scala 90:39]
  wire [24:0] _T_597; // @[Shift.scala 90:39]
  wire  _T_598; // @[Shift.scala 12:21]
  wire  _T_599; // @[Shift.scala 12:21]
  wire [1:0] _T_601; // @[Bitwise.scala 71:12]
  wire [26:0] _T_602; // @[Cat.scala 29:58]
  wire [26:0] _T_603; // @[Shift.scala 91:22]
  wire  _T_604; // @[Shift.scala 92:77]
  wire [25:0] _T_605; // @[Shift.scala 90:30]
  wire  _T_606; // @[Shift.scala 90:48]
  wire [25:0] _GEN_18; // @[Shift.scala 90:39]
  wire [25:0] _T_608; // @[Shift.scala 90:39]
  wire  _T_610; // @[Shift.scala 12:21]
  wire [26:0] _T_611; // @[Cat.scala 29:58]
  wire [26:0] _T_612; // @[Shift.scala 91:22]
  wire [26:0] _T_615; // @[Bitwise.scala 71:12]
  wire [26:0] smallerSig; // @[Shift.scala 39:10]
  wire [27:0] rawSumSig; // @[PositFMA.scala 118:34]
  wire  _T_616; // @[PositFMA.scala 119:42]
  wire  _T_617; // @[PositFMA.scala 119:46]
  wire  _T_618; // @[PositFMA.scala 119:79]
  wire  sumSign; // @[PositFMA.scala 119:63]
  wire [26:0] _T_620; // @[PositFMA.scala 120:50]
  wire [27:0] signSumSig; // @[Cat.scala 29:58]
  wire [26:0] _T_621; // @[PositFMA.scala 124:33]
  wire [26:0] _T_622; // @[PositFMA.scala 124:68]
  wire [26:0] sumXor; // @[PositFMA.scala 124:51]
  wire [15:0] _T_623; // @[LZD.scala 43:32]
  wire [7:0] _T_624; // @[LZD.scala 43:32]
  wire [3:0] _T_625; // @[LZD.scala 43:32]
  wire [1:0] _T_626; // @[LZD.scala 43:32]
  wire  _T_627; // @[LZD.scala 39:14]
  wire  _T_628; // @[LZD.scala 39:21]
  wire  _T_629; // @[LZD.scala 39:30]
  wire  _T_630; // @[LZD.scala 39:27]
  wire  _T_631; // @[LZD.scala 39:25]
  wire [1:0] _T_632; // @[Cat.scala 29:58]
  wire [1:0] _T_633; // @[LZD.scala 44:32]
  wire  _T_634; // @[LZD.scala 39:14]
  wire  _T_635; // @[LZD.scala 39:21]
  wire  _T_636; // @[LZD.scala 39:30]
  wire  _T_637; // @[LZD.scala 39:27]
  wire  _T_638; // @[LZD.scala 39:25]
  wire [1:0] _T_639; // @[Cat.scala 29:58]
  wire  _T_640; // @[Shift.scala 12:21]
  wire  _T_641; // @[Shift.scala 12:21]
  wire  _T_642; // @[LZD.scala 49:16]
  wire  _T_643; // @[LZD.scala 49:27]
  wire  _T_644; // @[LZD.scala 49:25]
  wire  _T_645; // @[LZD.scala 49:47]
  wire  _T_646; // @[LZD.scala 49:59]
  wire  _T_647; // @[LZD.scala 49:35]
  wire [2:0] _T_649; // @[Cat.scala 29:58]
  wire [3:0] _T_650; // @[LZD.scala 44:32]
  wire [1:0] _T_651; // @[LZD.scala 43:32]
  wire  _T_652; // @[LZD.scala 39:14]
  wire  _T_653; // @[LZD.scala 39:21]
  wire  _T_654; // @[LZD.scala 39:30]
  wire  _T_655; // @[LZD.scala 39:27]
  wire  _T_656; // @[LZD.scala 39:25]
  wire [1:0] _T_657; // @[Cat.scala 29:58]
  wire [1:0] _T_658; // @[LZD.scala 44:32]
  wire  _T_659; // @[LZD.scala 39:14]
  wire  _T_660; // @[LZD.scala 39:21]
  wire  _T_661; // @[LZD.scala 39:30]
  wire  _T_662; // @[LZD.scala 39:27]
  wire  _T_663; // @[LZD.scala 39:25]
  wire [1:0] _T_664; // @[Cat.scala 29:58]
  wire  _T_665; // @[Shift.scala 12:21]
  wire  _T_666; // @[Shift.scala 12:21]
  wire  _T_667; // @[LZD.scala 49:16]
  wire  _T_668; // @[LZD.scala 49:27]
  wire  _T_669; // @[LZD.scala 49:25]
  wire  _T_670; // @[LZD.scala 49:47]
  wire  _T_671; // @[LZD.scala 49:59]
  wire  _T_672; // @[LZD.scala 49:35]
  wire [2:0] _T_674; // @[Cat.scala 29:58]
  wire  _T_675; // @[Shift.scala 12:21]
  wire  _T_676; // @[Shift.scala 12:21]
  wire  _T_677; // @[LZD.scala 49:16]
  wire  _T_678; // @[LZD.scala 49:27]
  wire  _T_679; // @[LZD.scala 49:25]
  wire [1:0] _T_680; // @[LZD.scala 49:47]
  wire [1:0] _T_681; // @[LZD.scala 49:59]
  wire [1:0] _T_682; // @[LZD.scala 49:35]
  wire [3:0] _T_684; // @[Cat.scala 29:58]
  wire [7:0] _T_685; // @[LZD.scala 44:32]
  wire [3:0] _T_686; // @[LZD.scala 43:32]
  wire [1:0] _T_687; // @[LZD.scala 43:32]
  wire  _T_688; // @[LZD.scala 39:14]
  wire  _T_689; // @[LZD.scala 39:21]
  wire  _T_690; // @[LZD.scala 39:30]
  wire  _T_691; // @[LZD.scala 39:27]
  wire  _T_692; // @[LZD.scala 39:25]
  wire [1:0] _T_693; // @[Cat.scala 29:58]
  wire [1:0] _T_694; // @[LZD.scala 44:32]
  wire  _T_695; // @[LZD.scala 39:14]
  wire  _T_696; // @[LZD.scala 39:21]
  wire  _T_697; // @[LZD.scala 39:30]
  wire  _T_698; // @[LZD.scala 39:27]
  wire  _T_699; // @[LZD.scala 39:25]
  wire [1:0] _T_700; // @[Cat.scala 29:58]
  wire  _T_701; // @[Shift.scala 12:21]
  wire  _T_702; // @[Shift.scala 12:21]
  wire  _T_703; // @[LZD.scala 49:16]
  wire  _T_704; // @[LZD.scala 49:27]
  wire  _T_705; // @[LZD.scala 49:25]
  wire  _T_706; // @[LZD.scala 49:47]
  wire  _T_707; // @[LZD.scala 49:59]
  wire  _T_708; // @[LZD.scala 49:35]
  wire [2:0] _T_710; // @[Cat.scala 29:58]
  wire [3:0] _T_711; // @[LZD.scala 44:32]
  wire [1:0] _T_712; // @[LZD.scala 43:32]
  wire  _T_713; // @[LZD.scala 39:14]
  wire  _T_714; // @[LZD.scala 39:21]
  wire  _T_715; // @[LZD.scala 39:30]
  wire  _T_716; // @[LZD.scala 39:27]
  wire  _T_717; // @[LZD.scala 39:25]
  wire [1:0] _T_718; // @[Cat.scala 29:58]
  wire [1:0] _T_719; // @[LZD.scala 44:32]
  wire  _T_720; // @[LZD.scala 39:14]
  wire  _T_721; // @[LZD.scala 39:21]
  wire  _T_722; // @[LZD.scala 39:30]
  wire  _T_723; // @[LZD.scala 39:27]
  wire  _T_724; // @[LZD.scala 39:25]
  wire [1:0] _T_725; // @[Cat.scala 29:58]
  wire  _T_726; // @[Shift.scala 12:21]
  wire  _T_727; // @[Shift.scala 12:21]
  wire  _T_728; // @[LZD.scala 49:16]
  wire  _T_729; // @[LZD.scala 49:27]
  wire  _T_730; // @[LZD.scala 49:25]
  wire  _T_731; // @[LZD.scala 49:47]
  wire  _T_732; // @[LZD.scala 49:59]
  wire  _T_733; // @[LZD.scala 49:35]
  wire [2:0] _T_735; // @[Cat.scala 29:58]
  wire  _T_736; // @[Shift.scala 12:21]
  wire  _T_737; // @[Shift.scala 12:21]
  wire  _T_738; // @[LZD.scala 49:16]
  wire  _T_739; // @[LZD.scala 49:27]
  wire  _T_740; // @[LZD.scala 49:25]
  wire [1:0] _T_741; // @[LZD.scala 49:47]
  wire [1:0] _T_742; // @[LZD.scala 49:59]
  wire [1:0] _T_743; // @[LZD.scala 49:35]
  wire [3:0] _T_745; // @[Cat.scala 29:58]
  wire  _T_746; // @[Shift.scala 12:21]
  wire  _T_747; // @[Shift.scala 12:21]
  wire  _T_748; // @[LZD.scala 49:16]
  wire  _T_749; // @[LZD.scala 49:27]
  wire  _T_750; // @[LZD.scala 49:25]
  wire [2:0] _T_751; // @[LZD.scala 49:47]
  wire [2:0] _T_752; // @[LZD.scala 49:59]
  wire [2:0] _T_753; // @[LZD.scala 49:35]
  wire [4:0] _T_755; // @[Cat.scala 29:58]
  wire [10:0] _T_756; // @[LZD.scala 44:32]
  wire [7:0] _T_757; // @[LZD.scala 43:32]
  wire [3:0] _T_758; // @[LZD.scala 43:32]
  wire [1:0] _T_759; // @[LZD.scala 43:32]
  wire  _T_760; // @[LZD.scala 39:14]
  wire  _T_761; // @[LZD.scala 39:21]
  wire  _T_762; // @[LZD.scala 39:30]
  wire  _T_763; // @[LZD.scala 39:27]
  wire  _T_764; // @[LZD.scala 39:25]
  wire [1:0] _T_765; // @[Cat.scala 29:58]
  wire [1:0] _T_766; // @[LZD.scala 44:32]
  wire  _T_767; // @[LZD.scala 39:14]
  wire  _T_768; // @[LZD.scala 39:21]
  wire  _T_769; // @[LZD.scala 39:30]
  wire  _T_770; // @[LZD.scala 39:27]
  wire  _T_771; // @[LZD.scala 39:25]
  wire [1:0] _T_772; // @[Cat.scala 29:58]
  wire  _T_773; // @[Shift.scala 12:21]
  wire  _T_774; // @[Shift.scala 12:21]
  wire  _T_775; // @[LZD.scala 49:16]
  wire  _T_776; // @[LZD.scala 49:27]
  wire  _T_777; // @[LZD.scala 49:25]
  wire  _T_778; // @[LZD.scala 49:47]
  wire  _T_779; // @[LZD.scala 49:59]
  wire  _T_780; // @[LZD.scala 49:35]
  wire [2:0] _T_782; // @[Cat.scala 29:58]
  wire [3:0] _T_783; // @[LZD.scala 44:32]
  wire [1:0] _T_784; // @[LZD.scala 43:32]
  wire  _T_785; // @[LZD.scala 39:14]
  wire  _T_786; // @[LZD.scala 39:21]
  wire  _T_787; // @[LZD.scala 39:30]
  wire  _T_788; // @[LZD.scala 39:27]
  wire  _T_789; // @[LZD.scala 39:25]
  wire [1:0] _T_790; // @[Cat.scala 29:58]
  wire [1:0] _T_791; // @[LZD.scala 44:32]
  wire  _T_792; // @[LZD.scala 39:14]
  wire  _T_793; // @[LZD.scala 39:21]
  wire  _T_794; // @[LZD.scala 39:30]
  wire  _T_795; // @[LZD.scala 39:27]
  wire  _T_796; // @[LZD.scala 39:25]
  wire [1:0] _T_797; // @[Cat.scala 29:58]
  wire  _T_798; // @[Shift.scala 12:21]
  wire  _T_799; // @[Shift.scala 12:21]
  wire  _T_800; // @[LZD.scala 49:16]
  wire  _T_801; // @[LZD.scala 49:27]
  wire  _T_802; // @[LZD.scala 49:25]
  wire  _T_803; // @[LZD.scala 49:47]
  wire  _T_804; // @[LZD.scala 49:59]
  wire  _T_805; // @[LZD.scala 49:35]
  wire [2:0] _T_807; // @[Cat.scala 29:58]
  wire  _T_808; // @[Shift.scala 12:21]
  wire  _T_809; // @[Shift.scala 12:21]
  wire  _T_810; // @[LZD.scala 49:16]
  wire  _T_811; // @[LZD.scala 49:27]
  wire  _T_812; // @[LZD.scala 49:25]
  wire [1:0] _T_813; // @[LZD.scala 49:47]
  wire [1:0] _T_814; // @[LZD.scala 49:59]
  wire [1:0] _T_815; // @[LZD.scala 49:35]
  wire [3:0] _T_817; // @[Cat.scala 29:58]
  wire [2:0] _T_818; // @[LZD.scala 44:32]
  wire [1:0] _T_819; // @[LZD.scala 43:32]
  wire  _T_820; // @[LZD.scala 39:14]
  wire  _T_821; // @[LZD.scala 39:21]
  wire  _T_822; // @[LZD.scala 39:30]
  wire  _T_823; // @[LZD.scala 39:27]
  wire  _T_824; // @[LZD.scala 39:25]
  wire [1:0] _T_825; // @[Cat.scala 29:58]
  wire  _T_826; // @[LZD.scala 44:32]
  wire  _T_828; // @[Shift.scala 12:21]
  wire  _T_830; // @[LZD.scala 55:32]
  wire  _T_831; // @[LZD.scala 55:20]
  wire  _T_833; // @[Shift.scala 12:21]
  wire [2:0] _T_835; // @[Cat.scala 29:58]
  wire [2:0] _T_836; // @[LZD.scala 55:32]
  wire [2:0] _T_837; // @[LZD.scala 55:20]
  wire [3:0] _T_838; // @[Cat.scala 29:58]
  wire  _T_839; // @[Shift.scala 12:21]
  wire [3:0] _T_841; // @[LZD.scala 55:32]
  wire [3:0] _T_842; // @[LZD.scala 55:20]
  wire [4:0] sumLZD; // @[Cat.scala 29:58]
  wire [4:0] shiftValue; // @[PositFMA.scala 126:24]
  wire [25:0] _T_843; // @[PositFMA.scala 127:38]
  wire  _T_844; // @[Shift.scala 16:24]
  wire  _T_846; // @[Shift.scala 12:21]
  wire [9:0] _T_847; // @[Shift.scala 64:52]
  wire [25:0] _T_849; // @[Cat.scala 29:58]
  wire [25:0] _T_850; // @[Shift.scala 64:27]
  wire [3:0] _T_851; // @[Shift.scala 66:70]
  wire  _T_852; // @[Shift.scala 12:21]
  wire [17:0] _T_853; // @[Shift.scala 64:52]
  wire [25:0] _T_855; // @[Cat.scala 29:58]
  wire [25:0] _T_856; // @[Shift.scala 64:27]
  wire [2:0] _T_857; // @[Shift.scala 66:70]
  wire  _T_858; // @[Shift.scala 12:21]
  wire [21:0] _T_859; // @[Shift.scala 64:52]
  wire [25:0] _T_861; // @[Cat.scala 29:58]
  wire [25:0] _T_862; // @[Shift.scala 64:27]
  wire [1:0] _T_863; // @[Shift.scala 66:70]
  wire  _T_864; // @[Shift.scala 12:21]
  wire [23:0] _T_865; // @[Shift.scala 64:52]
  wire [25:0] _T_867; // @[Cat.scala 29:58]
  wire [25:0] _T_868; // @[Shift.scala 64:27]
  wire  _T_869; // @[Shift.scala 66:70]
  wire [24:0] _T_871; // @[Shift.scala 64:52]
  wire [25:0] _T_872; // @[Cat.scala 29:58]
  wire [25:0] _T_873; // @[Shift.scala 64:27]
  wire [25:0] normalFracTmp; // @[Shift.scala 16:10]
  wire [6:0] _T_875; // @[PositFMA.scala 130:36]
  wire [6:0] _T_876; // @[PositFMA.scala 130:36]
  wire [5:0] _T_877; // @[Cat.scala 29:58]
  wire [5:0] _T_878; // @[PositFMA.scala 130:61]
  wire [6:0] _GEN_19; // @[PositFMA.scala 130:42]
  wire [6:0] _T_880; // @[PositFMA.scala 130:42]
  wire [6:0] sumScale; // @[PositFMA.scala 130:42]
  wire [11:0] sumFrac; // @[PositFMA.scala 131:41]
  wire [13:0] grsTmp; // @[PositFMA.scala 134:41]
  wire [1:0] _T_881; // @[PositFMA.scala 137:40]
  wire [11:0] _T_882; // @[PositFMA.scala 137:56]
  wire  _T_883; // @[PositFMA.scala 137:60]
  wire  underflow; // @[PositFMA.scala 144:32]
  wire  overflow; // @[PositFMA.scala 145:32]
  wire  _T_884; // @[PositFMA.scala 154:32]
  wire  decF_isZero; // @[PositFMA.scala 154:20]
  wire [6:0] _T_886; // @[Mux.scala 87:16]
  wire [6:0] _T_887; // @[Mux.scala 87:16]
  wire [5:0] _GEN_20; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  wire [5:0] decF_scale; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  wire  _T_888; // @[convert.scala 46:61]
  wire  _T_889; // @[convert.scala 46:52]
  wire  _T_891; // @[convert.scala 46:42]
  wire [4:0] _T_892; // @[convert.scala 48:34]
  wire  _T_893; // @[convert.scala 49:36]
  wire [4:0] _T_895; // @[convert.scala 50:36]
  wire [4:0] _T_896; // @[convert.scala 50:36]
  wire [4:0] _T_897; // @[convert.scala 50:28]
  wire  _T_898; // @[convert.scala 51:31]
  wire  _T_899; // @[convert.scala 52:43]
  wire [17:0] _T_903; // @[Cat.scala 29:58]
  wire [4:0] _T_904; // @[Shift.scala 39:17]
  wire  _T_905; // @[Shift.scala 39:24]
  wire [1:0] _T_907; // @[Shift.scala 90:30]
  wire [15:0] _T_908; // @[Shift.scala 90:48]
  wire  _T_909; // @[Shift.scala 90:57]
  wire [1:0] _GEN_21; // @[Shift.scala 90:39]
  wire [1:0] _T_910; // @[Shift.scala 90:39]
  wire  _T_911; // @[Shift.scala 12:21]
  wire  _T_912; // @[Shift.scala 12:21]
  wire [15:0] _T_914; // @[Bitwise.scala 71:12]
  wire [17:0] _T_915; // @[Cat.scala 29:58]
  wire [17:0] _T_916; // @[Shift.scala 91:22]
  wire [3:0] _T_917; // @[Shift.scala 92:77]
  wire [9:0] _T_918; // @[Shift.scala 90:30]
  wire [7:0] _T_919; // @[Shift.scala 90:48]
  wire  _T_920; // @[Shift.scala 90:57]
  wire [9:0] _GEN_22; // @[Shift.scala 90:39]
  wire [9:0] _T_921; // @[Shift.scala 90:39]
  wire  _T_922; // @[Shift.scala 12:21]
  wire  _T_923; // @[Shift.scala 12:21]
  wire [7:0] _T_925; // @[Bitwise.scala 71:12]
  wire [17:0] _T_926; // @[Cat.scala 29:58]
  wire [17:0] _T_927; // @[Shift.scala 91:22]
  wire [2:0] _T_928; // @[Shift.scala 92:77]
  wire [13:0] _T_929; // @[Shift.scala 90:30]
  wire [3:0] _T_930; // @[Shift.scala 90:48]
  wire  _T_931; // @[Shift.scala 90:57]
  wire [13:0] _GEN_23; // @[Shift.scala 90:39]
  wire [13:0] _T_932; // @[Shift.scala 90:39]
  wire  _T_933; // @[Shift.scala 12:21]
  wire  _T_934; // @[Shift.scala 12:21]
  wire [3:0] _T_936; // @[Bitwise.scala 71:12]
  wire [17:0] _T_937; // @[Cat.scala 29:58]
  wire [17:0] _T_938; // @[Shift.scala 91:22]
  wire [1:0] _T_939; // @[Shift.scala 92:77]
  wire [15:0] _T_940; // @[Shift.scala 90:30]
  wire [1:0] _T_941; // @[Shift.scala 90:48]
  wire  _T_942; // @[Shift.scala 90:57]
  wire [15:0] _GEN_24; // @[Shift.scala 90:39]
  wire [15:0] _T_943; // @[Shift.scala 90:39]
  wire  _T_944; // @[Shift.scala 12:21]
  wire  _T_945; // @[Shift.scala 12:21]
  wire [1:0] _T_947; // @[Bitwise.scala 71:12]
  wire [17:0] _T_948; // @[Cat.scala 29:58]
  wire [17:0] _T_949; // @[Shift.scala 91:22]
  wire  _T_950; // @[Shift.scala 92:77]
  wire [16:0] _T_951; // @[Shift.scala 90:30]
  wire  _T_952; // @[Shift.scala 90:48]
  wire [16:0] _GEN_25; // @[Shift.scala 90:39]
  wire [16:0] _T_954; // @[Shift.scala 90:39]
  wire  _T_956; // @[Shift.scala 12:21]
  wire [17:0] _T_957; // @[Cat.scala 29:58]
  wire [17:0] _T_958; // @[Shift.scala 91:22]
  wire [17:0] _T_961; // @[Bitwise.scala 71:12]
  wire [17:0] _T_962; // @[Shift.scala 39:10]
  wire  _T_963; // @[convert.scala 55:31]
  wire  _T_964; // @[convert.scala 56:31]
  wire  _T_965; // @[convert.scala 57:31]
  wire  _T_966; // @[convert.scala 58:31]
  wire [14:0] _T_967; // @[convert.scala 59:69]
  wire  _T_968; // @[convert.scala 59:81]
  wire  _T_969; // @[convert.scala 59:50]
  wire  _T_971; // @[convert.scala 60:81]
  wire  _T_972; // @[convert.scala 61:44]
  wire  _T_973; // @[convert.scala 61:52]
  wire  _T_974; // @[convert.scala 61:36]
  wire  _T_975; // @[convert.scala 62:63]
  wire  _T_976; // @[convert.scala 62:103]
  wire  _T_977; // @[convert.scala 62:60]
  wire [14:0] _GEN_26; // @[convert.scala 63:56]
  wire [14:0] _T_980; // @[convert.scala 63:56]
  wire [15:0] _T_981; // @[Cat.scala 29:58]
  reg  _T_985; // @[Valid.scala 117:22]
  reg [31:0] _RAND_8;
  reg [15:0] _T_989; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  assign _T = io_fmaOp[1]; // @[PositFMA.scala 47:36]
  assign _T_2 = _T ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_3 = _T_2 ^ io_A; // @[PositFMA.scala 47:41]
  assign _GEN_10 = {{15'd0}, _T}; // @[PositFMA.scala 47:49]
  assign realA = _T_3 + _GEN_10; // @[PositFMA.scala 47:49]
  assign _T_6 = io_fmaOp[0]; // @[PositFMA.scala 48:36]
  assign _T_8 = _T_6 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_9 = _T_8 ^ io_C; // @[PositFMA.scala 48:41]
  assign _GEN_11 = {{15'd0}, _T_6}; // @[PositFMA.scala 48:49]
  assign realC = _T_9 + _GEN_11; // @[PositFMA.scala 48:49]
  assign _T_13 = realA[15]; // @[convert.scala 18:24]
  assign _T_14 = realA[14]; // @[convert.scala 18:40]
  assign _T_15 = _T_13 ^ _T_14; // @[convert.scala 18:36]
  assign _T_16 = realA[14:1]; // @[convert.scala 19:24]
  assign _T_17 = realA[13:0]; // @[convert.scala 19:43]
  assign _T_18 = _T_16 ^ _T_17; // @[convert.scala 19:39]
  assign _T_19 = _T_18[13:6]; // @[LZD.scala 43:32]
  assign _T_20 = _T_19[7:4]; // @[LZD.scala 43:32]
  assign _T_21 = _T_20[3:2]; // @[LZD.scala 43:32]
  assign _T_22 = _T_21 != 2'h0; // @[LZD.scala 39:14]
  assign _T_23 = _T_21[1]; // @[LZD.scala 39:21]
  assign _T_24 = _T_21[0]; // @[LZD.scala 39:30]
  assign _T_25 = ~ _T_24; // @[LZD.scala 39:27]
  assign _T_26 = _T_23 | _T_25; // @[LZD.scala 39:25]
  assign _T_27 = {_T_22,_T_26}; // @[Cat.scala 29:58]
  assign _T_28 = _T_20[1:0]; // @[LZD.scala 44:32]
  assign _T_29 = _T_28 != 2'h0; // @[LZD.scala 39:14]
  assign _T_30 = _T_28[1]; // @[LZD.scala 39:21]
  assign _T_31 = _T_28[0]; // @[LZD.scala 39:30]
  assign _T_32 = ~ _T_31; // @[LZD.scala 39:27]
  assign _T_33 = _T_30 | _T_32; // @[LZD.scala 39:25]
  assign _T_34 = {_T_29,_T_33}; // @[Cat.scala 29:58]
  assign _T_35 = _T_27[1]; // @[Shift.scala 12:21]
  assign _T_36 = _T_34[1]; // @[Shift.scala 12:21]
  assign _T_37 = _T_35 | _T_36; // @[LZD.scala 49:16]
  assign _T_38 = ~ _T_36; // @[LZD.scala 49:27]
  assign _T_39 = _T_35 | _T_38; // @[LZD.scala 49:25]
  assign _T_40 = _T_27[0:0]; // @[LZD.scala 49:47]
  assign _T_41 = _T_34[0:0]; // @[LZD.scala 49:59]
  assign _T_42 = _T_35 ? _T_40 : _T_41; // @[LZD.scala 49:35]
  assign _T_44 = {_T_37,_T_39,_T_42}; // @[Cat.scala 29:58]
  assign _T_45 = _T_19[3:0]; // @[LZD.scala 44:32]
  assign _T_46 = _T_45[3:2]; // @[LZD.scala 43:32]
  assign _T_47 = _T_46 != 2'h0; // @[LZD.scala 39:14]
  assign _T_48 = _T_46[1]; // @[LZD.scala 39:21]
  assign _T_49 = _T_46[0]; // @[LZD.scala 39:30]
  assign _T_50 = ~ _T_49; // @[LZD.scala 39:27]
  assign _T_51 = _T_48 | _T_50; // @[LZD.scala 39:25]
  assign _T_52 = {_T_47,_T_51}; // @[Cat.scala 29:58]
  assign _T_53 = _T_45[1:0]; // @[LZD.scala 44:32]
  assign _T_54 = _T_53 != 2'h0; // @[LZD.scala 39:14]
  assign _T_55 = _T_53[1]; // @[LZD.scala 39:21]
  assign _T_56 = _T_53[0]; // @[LZD.scala 39:30]
  assign _T_57 = ~ _T_56; // @[LZD.scala 39:27]
  assign _T_58 = _T_55 | _T_57; // @[LZD.scala 39:25]
  assign _T_59 = {_T_54,_T_58}; // @[Cat.scala 29:58]
  assign _T_60 = _T_52[1]; // @[Shift.scala 12:21]
  assign _T_61 = _T_59[1]; // @[Shift.scala 12:21]
  assign _T_62 = _T_60 | _T_61; // @[LZD.scala 49:16]
  assign _T_63 = ~ _T_61; // @[LZD.scala 49:27]
  assign _T_64 = _T_60 | _T_63; // @[LZD.scala 49:25]
  assign _T_65 = _T_52[0:0]; // @[LZD.scala 49:47]
  assign _T_66 = _T_59[0:0]; // @[LZD.scala 49:59]
  assign _T_67 = _T_60 ? _T_65 : _T_66; // @[LZD.scala 49:35]
  assign _T_69 = {_T_62,_T_64,_T_67}; // @[Cat.scala 29:58]
  assign _T_70 = _T_44[2]; // @[Shift.scala 12:21]
  assign _T_71 = _T_69[2]; // @[Shift.scala 12:21]
  assign _T_72 = _T_70 | _T_71; // @[LZD.scala 49:16]
  assign _T_73 = ~ _T_71; // @[LZD.scala 49:27]
  assign _T_74 = _T_70 | _T_73; // @[LZD.scala 49:25]
  assign _T_75 = _T_44[1:0]; // @[LZD.scala 49:47]
  assign _T_76 = _T_69[1:0]; // @[LZD.scala 49:59]
  assign _T_77 = _T_70 ? _T_75 : _T_76; // @[LZD.scala 49:35]
  assign _T_79 = {_T_72,_T_74,_T_77}; // @[Cat.scala 29:58]
  assign _T_80 = _T_18[5:0]; // @[LZD.scala 44:32]
  assign _T_81 = _T_80[5:2]; // @[LZD.scala 43:32]
  assign _T_82 = _T_81[3:2]; // @[LZD.scala 43:32]
  assign _T_83 = _T_82 != 2'h0; // @[LZD.scala 39:14]
  assign _T_84 = _T_82[1]; // @[LZD.scala 39:21]
  assign _T_85 = _T_82[0]; // @[LZD.scala 39:30]
  assign _T_86 = ~ _T_85; // @[LZD.scala 39:27]
  assign _T_87 = _T_84 | _T_86; // @[LZD.scala 39:25]
  assign _T_88 = {_T_83,_T_87}; // @[Cat.scala 29:58]
  assign _T_89 = _T_81[1:0]; // @[LZD.scala 44:32]
  assign _T_90 = _T_89 != 2'h0; // @[LZD.scala 39:14]
  assign _T_91 = _T_89[1]; // @[LZD.scala 39:21]
  assign _T_92 = _T_89[0]; // @[LZD.scala 39:30]
  assign _T_93 = ~ _T_92; // @[LZD.scala 39:27]
  assign _T_94 = _T_91 | _T_93; // @[LZD.scala 39:25]
  assign _T_95 = {_T_90,_T_94}; // @[Cat.scala 29:58]
  assign _T_96 = _T_88[1]; // @[Shift.scala 12:21]
  assign _T_97 = _T_95[1]; // @[Shift.scala 12:21]
  assign _T_98 = _T_96 | _T_97; // @[LZD.scala 49:16]
  assign _T_99 = ~ _T_97; // @[LZD.scala 49:27]
  assign _T_100 = _T_96 | _T_99; // @[LZD.scala 49:25]
  assign _T_101 = _T_88[0:0]; // @[LZD.scala 49:47]
  assign _T_102 = _T_95[0:0]; // @[LZD.scala 49:59]
  assign _T_103 = _T_96 ? _T_101 : _T_102; // @[LZD.scala 49:35]
  assign _T_105 = {_T_98,_T_100,_T_103}; // @[Cat.scala 29:58]
  assign _T_106 = _T_80[1:0]; // @[LZD.scala 44:32]
  assign _T_107 = _T_106 != 2'h0; // @[LZD.scala 39:14]
  assign _T_108 = _T_106[1]; // @[LZD.scala 39:21]
  assign _T_109 = _T_106[0]; // @[LZD.scala 39:30]
  assign _T_110 = ~ _T_109; // @[LZD.scala 39:27]
  assign _T_111 = _T_108 | _T_110; // @[LZD.scala 39:25]
  assign _T_112 = {_T_107,_T_111}; // @[Cat.scala 29:58]
  assign _T_113 = _T_105[2]; // @[Shift.scala 12:21]
  assign _T_115 = _T_105[1:0]; // @[LZD.scala 55:32]
  assign _T_116 = _T_113 ? _T_115 : _T_112; // @[LZD.scala 55:20]
  assign _T_117 = {_T_113,_T_116}; // @[Cat.scala 29:58]
  assign _T_118 = _T_79[3]; // @[Shift.scala 12:21]
  assign _T_120 = _T_79[2:0]; // @[LZD.scala 55:32]
  assign _T_121 = _T_118 ? _T_120 : _T_117; // @[LZD.scala 55:20]
  assign _T_122 = {_T_118,_T_121}; // @[Cat.scala 29:58]
  assign _T_123 = ~ _T_122; // @[convert.scala 21:22]
  assign _T_124 = realA[12:0]; // @[convert.scala 22:36]
  assign _T_125 = _T_123 < 4'hd; // @[Shift.scala 16:24]
  assign _T_127 = _T_123[3]; // @[Shift.scala 12:21]
  assign _T_128 = _T_124[4:0]; // @[Shift.scala 64:52]
  assign _T_130 = {_T_128,8'h0}; // @[Cat.scala 29:58]
  assign _T_131 = _T_127 ? _T_130 : _T_124; // @[Shift.scala 64:27]
  assign _T_132 = _T_123[2:0]; // @[Shift.scala 66:70]
  assign _T_133 = _T_132[2]; // @[Shift.scala 12:21]
  assign _T_134 = _T_131[8:0]; // @[Shift.scala 64:52]
  assign _T_136 = {_T_134,4'h0}; // @[Cat.scala 29:58]
  assign _T_137 = _T_133 ? _T_136 : _T_131; // @[Shift.scala 64:27]
  assign _T_138 = _T_132[1:0]; // @[Shift.scala 66:70]
  assign _T_139 = _T_138[1]; // @[Shift.scala 12:21]
  assign _T_140 = _T_137[10:0]; // @[Shift.scala 64:52]
  assign _T_142 = {_T_140,2'h0}; // @[Cat.scala 29:58]
  assign _T_143 = _T_139 ? _T_142 : _T_137; // @[Shift.scala 64:27]
  assign _T_144 = _T_138[0:0]; // @[Shift.scala 66:70]
  assign _T_146 = _T_143[11:0]; // @[Shift.scala 64:52]
  assign _T_147 = {_T_146,1'h0}; // @[Cat.scala 29:58]
  assign _T_148 = _T_144 ? _T_147 : _T_143; // @[Shift.scala 64:27]
  assign _T_149 = _T_125 ? _T_148 : 13'h0; // @[Shift.scala 16:10]
  assign _T_150 = _T_149[12:12]; // @[convert.scala 23:34]
  assign decA_fraction = _T_149[11:0]; // @[convert.scala 24:34]
  assign _T_152 = _T_15 == 1'h0; // @[convert.scala 25:26]
  assign _T_154 = _T_15 ? _T_123 : _T_122; // @[convert.scala 25:42]
  assign _T_157 = ~ _T_150; // @[convert.scala 26:67]
  assign _T_158 = _T_13 ? _T_157 : _T_150; // @[convert.scala 26:51]
  assign _T_159 = {_T_152,_T_154,_T_158}; // @[Cat.scala 29:58]
  assign _T_161 = realA[14:0]; // @[convert.scala 29:56]
  assign _T_162 = _T_161 != 15'h0; // @[convert.scala 29:60]
  assign _T_163 = ~ _T_162; // @[convert.scala 29:41]
  assign decA_isNaR = _T_13 & _T_163; // @[convert.scala 29:39]
  assign _T_166 = _T_13 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_166 & _T_163; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_159); // @[convert.scala 32:24]
  assign _T_175 = io_B[15]; // @[convert.scala 18:24]
  assign _T_176 = io_B[14]; // @[convert.scala 18:40]
  assign _T_177 = _T_175 ^ _T_176; // @[convert.scala 18:36]
  assign _T_178 = io_B[14:1]; // @[convert.scala 19:24]
  assign _T_179 = io_B[13:0]; // @[convert.scala 19:43]
  assign _T_180 = _T_178 ^ _T_179; // @[convert.scala 19:39]
  assign _T_181 = _T_180[13:6]; // @[LZD.scala 43:32]
  assign _T_182 = _T_181[7:4]; // @[LZD.scala 43:32]
  assign _T_183 = _T_182[3:2]; // @[LZD.scala 43:32]
  assign _T_184 = _T_183 != 2'h0; // @[LZD.scala 39:14]
  assign _T_185 = _T_183[1]; // @[LZD.scala 39:21]
  assign _T_186 = _T_183[0]; // @[LZD.scala 39:30]
  assign _T_187 = ~ _T_186; // @[LZD.scala 39:27]
  assign _T_188 = _T_185 | _T_187; // @[LZD.scala 39:25]
  assign _T_189 = {_T_184,_T_188}; // @[Cat.scala 29:58]
  assign _T_190 = _T_182[1:0]; // @[LZD.scala 44:32]
  assign _T_191 = _T_190 != 2'h0; // @[LZD.scala 39:14]
  assign _T_192 = _T_190[1]; // @[LZD.scala 39:21]
  assign _T_193 = _T_190[0]; // @[LZD.scala 39:30]
  assign _T_194 = ~ _T_193; // @[LZD.scala 39:27]
  assign _T_195 = _T_192 | _T_194; // @[LZD.scala 39:25]
  assign _T_196 = {_T_191,_T_195}; // @[Cat.scala 29:58]
  assign _T_197 = _T_189[1]; // @[Shift.scala 12:21]
  assign _T_198 = _T_196[1]; // @[Shift.scala 12:21]
  assign _T_199 = _T_197 | _T_198; // @[LZD.scala 49:16]
  assign _T_200 = ~ _T_198; // @[LZD.scala 49:27]
  assign _T_201 = _T_197 | _T_200; // @[LZD.scala 49:25]
  assign _T_202 = _T_189[0:0]; // @[LZD.scala 49:47]
  assign _T_203 = _T_196[0:0]; // @[LZD.scala 49:59]
  assign _T_204 = _T_197 ? _T_202 : _T_203; // @[LZD.scala 49:35]
  assign _T_206 = {_T_199,_T_201,_T_204}; // @[Cat.scala 29:58]
  assign _T_207 = _T_181[3:0]; // @[LZD.scala 44:32]
  assign _T_208 = _T_207[3:2]; // @[LZD.scala 43:32]
  assign _T_209 = _T_208 != 2'h0; // @[LZD.scala 39:14]
  assign _T_210 = _T_208[1]; // @[LZD.scala 39:21]
  assign _T_211 = _T_208[0]; // @[LZD.scala 39:30]
  assign _T_212 = ~ _T_211; // @[LZD.scala 39:27]
  assign _T_213 = _T_210 | _T_212; // @[LZD.scala 39:25]
  assign _T_214 = {_T_209,_T_213}; // @[Cat.scala 29:58]
  assign _T_215 = _T_207[1:0]; // @[LZD.scala 44:32]
  assign _T_216 = _T_215 != 2'h0; // @[LZD.scala 39:14]
  assign _T_217 = _T_215[1]; // @[LZD.scala 39:21]
  assign _T_218 = _T_215[0]; // @[LZD.scala 39:30]
  assign _T_219 = ~ _T_218; // @[LZD.scala 39:27]
  assign _T_220 = _T_217 | _T_219; // @[LZD.scala 39:25]
  assign _T_221 = {_T_216,_T_220}; // @[Cat.scala 29:58]
  assign _T_222 = _T_214[1]; // @[Shift.scala 12:21]
  assign _T_223 = _T_221[1]; // @[Shift.scala 12:21]
  assign _T_224 = _T_222 | _T_223; // @[LZD.scala 49:16]
  assign _T_225 = ~ _T_223; // @[LZD.scala 49:27]
  assign _T_226 = _T_222 | _T_225; // @[LZD.scala 49:25]
  assign _T_227 = _T_214[0:0]; // @[LZD.scala 49:47]
  assign _T_228 = _T_221[0:0]; // @[LZD.scala 49:59]
  assign _T_229 = _T_222 ? _T_227 : _T_228; // @[LZD.scala 49:35]
  assign _T_231 = {_T_224,_T_226,_T_229}; // @[Cat.scala 29:58]
  assign _T_232 = _T_206[2]; // @[Shift.scala 12:21]
  assign _T_233 = _T_231[2]; // @[Shift.scala 12:21]
  assign _T_234 = _T_232 | _T_233; // @[LZD.scala 49:16]
  assign _T_235 = ~ _T_233; // @[LZD.scala 49:27]
  assign _T_236 = _T_232 | _T_235; // @[LZD.scala 49:25]
  assign _T_237 = _T_206[1:0]; // @[LZD.scala 49:47]
  assign _T_238 = _T_231[1:0]; // @[LZD.scala 49:59]
  assign _T_239 = _T_232 ? _T_237 : _T_238; // @[LZD.scala 49:35]
  assign _T_241 = {_T_234,_T_236,_T_239}; // @[Cat.scala 29:58]
  assign _T_242 = _T_180[5:0]; // @[LZD.scala 44:32]
  assign _T_243 = _T_242[5:2]; // @[LZD.scala 43:32]
  assign _T_244 = _T_243[3:2]; // @[LZD.scala 43:32]
  assign _T_245 = _T_244 != 2'h0; // @[LZD.scala 39:14]
  assign _T_246 = _T_244[1]; // @[LZD.scala 39:21]
  assign _T_247 = _T_244[0]; // @[LZD.scala 39:30]
  assign _T_248 = ~ _T_247; // @[LZD.scala 39:27]
  assign _T_249 = _T_246 | _T_248; // @[LZD.scala 39:25]
  assign _T_250 = {_T_245,_T_249}; // @[Cat.scala 29:58]
  assign _T_251 = _T_243[1:0]; // @[LZD.scala 44:32]
  assign _T_252 = _T_251 != 2'h0; // @[LZD.scala 39:14]
  assign _T_253 = _T_251[1]; // @[LZD.scala 39:21]
  assign _T_254 = _T_251[0]; // @[LZD.scala 39:30]
  assign _T_255 = ~ _T_254; // @[LZD.scala 39:27]
  assign _T_256 = _T_253 | _T_255; // @[LZD.scala 39:25]
  assign _T_257 = {_T_252,_T_256}; // @[Cat.scala 29:58]
  assign _T_258 = _T_250[1]; // @[Shift.scala 12:21]
  assign _T_259 = _T_257[1]; // @[Shift.scala 12:21]
  assign _T_260 = _T_258 | _T_259; // @[LZD.scala 49:16]
  assign _T_261 = ~ _T_259; // @[LZD.scala 49:27]
  assign _T_262 = _T_258 | _T_261; // @[LZD.scala 49:25]
  assign _T_263 = _T_250[0:0]; // @[LZD.scala 49:47]
  assign _T_264 = _T_257[0:0]; // @[LZD.scala 49:59]
  assign _T_265 = _T_258 ? _T_263 : _T_264; // @[LZD.scala 49:35]
  assign _T_267 = {_T_260,_T_262,_T_265}; // @[Cat.scala 29:58]
  assign _T_268 = _T_242[1:0]; // @[LZD.scala 44:32]
  assign _T_269 = _T_268 != 2'h0; // @[LZD.scala 39:14]
  assign _T_270 = _T_268[1]; // @[LZD.scala 39:21]
  assign _T_271 = _T_268[0]; // @[LZD.scala 39:30]
  assign _T_272 = ~ _T_271; // @[LZD.scala 39:27]
  assign _T_273 = _T_270 | _T_272; // @[LZD.scala 39:25]
  assign _T_274 = {_T_269,_T_273}; // @[Cat.scala 29:58]
  assign _T_275 = _T_267[2]; // @[Shift.scala 12:21]
  assign _T_277 = _T_267[1:0]; // @[LZD.scala 55:32]
  assign _T_278 = _T_275 ? _T_277 : _T_274; // @[LZD.scala 55:20]
  assign _T_279 = {_T_275,_T_278}; // @[Cat.scala 29:58]
  assign _T_280 = _T_241[3]; // @[Shift.scala 12:21]
  assign _T_282 = _T_241[2:0]; // @[LZD.scala 55:32]
  assign _T_283 = _T_280 ? _T_282 : _T_279; // @[LZD.scala 55:20]
  assign _T_284 = {_T_280,_T_283}; // @[Cat.scala 29:58]
  assign _T_285 = ~ _T_284; // @[convert.scala 21:22]
  assign _T_286 = io_B[12:0]; // @[convert.scala 22:36]
  assign _T_287 = _T_285 < 4'hd; // @[Shift.scala 16:24]
  assign _T_289 = _T_285[3]; // @[Shift.scala 12:21]
  assign _T_290 = _T_286[4:0]; // @[Shift.scala 64:52]
  assign _T_292 = {_T_290,8'h0}; // @[Cat.scala 29:58]
  assign _T_293 = _T_289 ? _T_292 : _T_286; // @[Shift.scala 64:27]
  assign _T_294 = _T_285[2:0]; // @[Shift.scala 66:70]
  assign _T_295 = _T_294[2]; // @[Shift.scala 12:21]
  assign _T_296 = _T_293[8:0]; // @[Shift.scala 64:52]
  assign _T_298 = {_T_296,4'h0}; // @[Cat.scala 29:58]
  assign _T_299 = _T_295 ? _T_298 : _T_293; // @[Shift.scala 64:27]
  assign _T_300 = _T_294[1:0]; // @[Shift.scala 66:70]
  assign _T_301 = _T_300[1]; // @[Shift.scala 12:21]
  assign _T_302 = _T_299[10:0]; // @[Shift.scala 64:52]
  assign _T_304 = {_T_302,2'h0}; // @[Cat.scala 29:58]
  assign _T_305 = _T_301 ? _T_304 : _T_299; // @[Shift.scala 64:27]
  assign _T_306 = _T_300[0:0]; // @[Shift.scala 66:70]
  assign _T_308 = _T_305[11:0]; // @[Shift.scala 64:52]
  assign _T_309 = {_T_308,1'h0}; // @[Cat.scala 29:58]
  assign _T_310 = _T_306 ? _T_309 : _T_305; // @[Shift.scala 64:27]
  assign _T_311 = _T_287 ? _T_310 : 13'h0; // @[Shift.scala 16:10]
  assign _T_312 = _T_311[12:12]; // @[convert.scala 23:34]
  assign decB_fraction = _T_311[11:0]; // @[convert.scala 24:34]
  assign _T_314 = _T_177 == 1'h0; // @[convert.scala 25:26]
  assign _T_316 = _T_177 ? _T_285 : _T_284; // @[convert.scala 25:42]
  assign _T_319 = ~ _T_312; // @[convert.scala 26:67]
  assign _T_320 = _T_175 ? _T_319 : _T_312; // @[convert.scala 26:51]
  assign _T_321 = {_T_314,_T_316,_T_320}; // @[Cat.scala 29:58]
  assign _T_323 = io_B[14:0]; // @[convert.scala 29:56]
  assign _T_324 = _T_323 != 15'h0; // @[convert.scala 29:60]
  assign _T_325 = ~ _T_324; // @[convert.scala 29:41]
  assign decB_isNaR = _T_175 & _T_325; // @[convert.scala 29:39]
  assign _T_328 = _T_175 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_328 & _T_325; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_321); // @[convert.scala 32:24]
  assign _T_337 = realC[15]; // @[convert.scala 18:24]
  assign _T_338 = realC[14]; // @[convert.scala 18:40]
  assign _T_339 = _T_337 ^ _T_338; // @[convert.scala 18:36]
  assign _T_340 = realC[14:1]; // @[convert.scala 19:24]
  assign _T_341 = realC[13:0]; // @[convert.scala 19:43]
  assign _T_342 = _T_340 ^ _T_341; // @[convert.scala 19:39]
  assign _T_343 = _T_342[13:6]; // @[LZD.scala 43:32]
  assign _T_344 = _T_343[7:4]; // @[LZD.scala 43:32]
  assign _T_345 = _T_344[3:2]; // @[LZD.scala 43:32]
  assign _T_346 = _T_345 != 2'h0; // @[LZD.scala 39:14]
  assign _T_347 = _T_345[1]; // @[LZD.scala 39:21]
  assign _T_348 = _T_345[0]; // @[LZD.scala 39:30]
  assign _T_349 = ~ _T_348; // @[LZD.scala 39:27]
  assign _T_350 = _T_347 | _T_349; // @[LZD.scala 39:25]
  assign _T_351 = {_T_346,_T_350}; // @[Cat.scala 29:58]
  assign _T_352 = _T_344[1:0]; // @[LZD.scala 44:32]
  assign _T_353 = _T_352 != 2'h0; // @[LZD.scala 39:14]
  assign _T_354 = _T_352[1]; // @[LZD.scala 39:21]
  assign _T_355 = _T_352[0]; // @[LZD.scala 39:30]
  assign _T_356 = ~ _T_355; // @[LZD.scala 39:27]
  assign _T_357 = _T_354 | _T_356; // @[LZD.scala 39:25]
  assign _T_358 = {_T_353,_T_357}; // @[Cat.scala 29:58]
  assign _T_359 = _T_351[1]; // @[Shift.scala 12:21]
  assign _T_360 = _T_358[1]; // @[Shift.scala 12:21]
  assign _T_361 = _T_359 | _T_360; // @[LZD.scala 49:16]
  assign _T_362 = ~ _T_360; // @[LZD.scala 49:27]
  assign _T_363 = _T_359 | _T_362; // @[LZD.scala 49:25]
  assign _T_364 = _T_351[0:0]; // @[LZD.scala 49:47]
  assign _T_365 = _T_358[0:0]; // @[LZD.scala 49:59]
  assign _T_366 = _T_359 ? _T_364 : _T_365; // @[LZD.scala 49:35]
  assign _T_368 = {_T_361,_T_363,_T_366}; // @[Cat.scala 29:58]
  assign _T_369 = _T_343[3:0]; // @[LZD.scala 44:32]
  assign _T_370 = _T_369[3:2]; // @[LZD.scala 43:32]
  assign _T_371 = _T_370 != 2'h0; // @[LZD.scala 39:14]
  assign _T_372 = _T_370[1]; // @[LZD.scala 39:21]
  assign _T_373 = _T_370[0]; // @[LZD.scala 39:30]
  assign _T_374 = ~ _T_373; // @[LZD.scala 39:27]
  assign _T_375 = _T_372 | _T_374; // @[LZD.scala 39:25]
  assign _T_376 = {_T_371,_T_375}; // @[Cat.scala 29:58]
  assign _T_377 = _T_369[1:0]; // @[LZD.scala 44:32]
  assign _T_378 = _T_377 != 2'h0; // @[LZD.scala 39:14]
  assign _T_379 = _T_377[1]; // @[LZD.scala 39:21]
  assign _T_380 = _T_377[0]; // @[LZD.scala 39:30]
  assign _T_381 = ~ _T_380; // @[LZD.scala 39:27]
  assign _T_382 = _T_379 | _T_381; // @[LZD.scala 39:25]
  assign _T_383 = {_T_378,_T_382}; // @[Cat.scala 29:58]
  assign _T_384 = _T_376[1]; // @[Shift.scala 12:21]
  assign _T_385 = _T_383[1]; // @[Shift.scala 12:21]
  assign _T_386 = _T_384 | _T_385; // @[LZD.scala 49:16]
  assign _T_387 = ~ _T_385; // @[LZD.scala 49:27]
  assign _T_388 = _T_384 | _T_387; // @[LZD.scala 49:25]
  assign _T_389 = _T_376[0:0]; // @[LZD.scala 49:47]
  assign _T_390 = _T_383[0:0]; // @[LZD.scala 49:59]
  assign _T_391 = _T_384 ? _T_389 : _T_390; // @[LZD.scala 49:35]
  assign _T_393 = {_T_386,_T_388,_T_391}; // @[Cat.scala 29:58]
  assign _T_394 = _T_368[2]; // @[Shift.scala 12:21]
  assign _T_395 = _T_393[2]; // @[Shift.scala 12:21]
  assign _T_396 = _T_394 | _T_395; // @[LZD.scala 49:16]
  assign _T_397 = ~ _T_395; // @[LZD.scala 49:27]
  assign _T_398 = _T_394 | _T_397; // @[LZD.scala 49:25]
  assign _T_399 = _T_368[1:0]; // @[LZD.scala 49:47]
  assign _T_400 = _T_393[1:0]; // @[LZD.scala 49:59]
  assign _T_401 = _T_394 ? _T_399 : _T_400; // @[LZD.scala 49:35]
  assign _T_403 = {_T_396,_T_398,_T_401}; // @[Cat.scala 29:58]
  assign _T_404 = _T_342[5:0]; // @[LZD.scala 44:32]
  assign _T_405 = _T_404[5:2]; // @[LZD.scala 43:32]
  assign _T_406 = _T_405[3:2]; // @[LZD.scala 43:32]
  assign _T_407 = _T_406 != 2'h0; // @[LZD.scala 39:14]
  assign _T_408 = _T_406[1]; // @[LZD.scala 39:21]
  assign _T_409 = _T_406[0]; // @[LZD.scala 39:30]
  assign _T_410 = ~ _T_409; // @[LZD.scala 39:27]
  assign _T_411 = _T_408 | _T_410; // @[LZD.scala 39:25]
  assign _T_412 = {_T_407,_T_411}; // @[Cat.scala 29:58]
  assign _T_413 = _T_405[1:0]; // @[LZD.scala 44:32]
  assign _T_414 = _T_413 != 2'h0; // @[LZD.scala 39:14]
  assign _T_415 = _T_413[1]; // @[LZD.scala 39:21]
  assign _T_416 = _T_413[0]; // @[LZD.scala 39:30]
  assign _T_417 = ~ _T_416; // @[LZD.scala 39:27]
  assign _T_418 = _T_415 | _T_417; // @[LZD.scala 39:25]
  assign _T_419 = {_T_414,_T_418}; // @[Cat.scala 29:58]
  assign _T_420 = _T_412[1]; // @[Shift.scala 12:21]
  assign _T_421 = _T_419[1]; // @[Shift.scala 12:21]
  assign _T_422 = _T_420 | _T_421; // @[LZD.scala 49:16]
  assign _T_423 = ~ _T_421; // @[LZD.scala 49:27]
  assign _T_424 = _T_420 | _T_423; // @[LZD.scala 49:25]
  assign _T_425 = _T_412[0:0]; // @[LZD.scala 49:47]
  assign _T_426 = _T_419[0:0]; // @[LZD.scala 49:59]
  assign _T_427 = _T_420 ? _T_425 : _T_426; // @[LZD.scala 49:35]
  assign _T_429 = {_T_422,_T_424,_T_427}; // @[Cat.scala 29:58]
  assign _T_430 = _T_404[1:0]; // @[LZD.scala 44:32]
  assign _T_431 = _T_430 != 2'h0; // @[LZD.scala 39:14]
  assign _T_432 = _T_430[1]; // @[LZD.scala 39:21]
  assign _T_433 = _T_430[0]; // @[LZD.scala 39:30]
  assign _T_434 = ~ _T_433; // @[LZD.scala 39:27]
  assign _T_435 = _T_432 | _T_434; // @[LZD.scala 39:25]
  assign _T_436 = {_T_431,_T_435}; // @[Cat.scala 29:58]
  assign _T_437 = _T_429[2]; // @[Shift.scala 12:21]
  assign _T_439 = _T_429[1:0]; // @[LZD.scala 55:32]
  assign _T_440 = _T_437 ? _T_439 : _T_436; // @[LZD.scala 55:20]
  assign _T_441 = {_T_437,_T_440}; // @[Cat.scala 29:58]
  assign _T_442 = _T_403[3]; // @[Shift.scala 12:21]
  assign _T_444 = _T_403[2:0]; // @[LZD.scala 55:32]
  assign _T_445 = _T_442 ? _T_444 : _T_441; // @[LZD.scala 55:20]
  assign _T_446 = {_T_442,_T_445}; // @[Cat.scala 29:58]
  assign _T_447 = ~ _T_446; // @[convert.scala 21:22]
  assign _T_448 = realC[12:0]; // @[convert.scala 22:36]
  assign _T_449 = _T_447 < 4'hd; // @[Shift.scala 16:24]
  assign _T_451 = _T_447[3]; // @[Shift.scala 12:21]
  assign _T_452 = _T_448[4:0]; // @[Shift.scala 64:52]
  assign _T_454 = {_T_452,8'h0}; // @[Cat.scala 29:58]
  assign _T_455 = _T_451 ? _T_454 : _T_448; // @[Shift.scala 64:27]
  assign _T_456 = _T_447[2:0]; // @[Shift.scala 66:70]
  assign _T_457 = _T_456[2]; // @[Shift.scala 12:21]
  assign _T_458 = _T_455[8:0]; // @[Shift.scala 64:52]
  assign _T_460 = {_T_458,4'h0}; // @[Cat.scala 29:58]
  assign _T_461 = _T_457 ? _T_460 : _T_455; // @[Shift.scala 64:27]
  assign _T_462 = _T_456[1:0]; // @[Shift.scala 66:70]
  assign _T_463 = _T_462[1]; // @[Shift.scala 12:21]
  assign _T_464 = _T_461[10:0]; // @[Shift.scala 64:52]
  assign _T_466 = {_T_464,2'h0}; // @[Cat.scala 29:58]
  assign _T_467 = _T_463 ? _T_466 : _T_461; // @[Shift.scala 64:27]
  assign _T_468 = _T_462[0:0]; // @[Shift.scala 66:70]
  assign _T_470 = _T_467[11:0]; // @[Shift.scala 64:52]
  assign _T_471 = {_T_470,1'h0}; // @[Cat.scala 29:58]
  assign _T_472 = _T_468 ? _T_471 : _T_467; // @[Shift.scala 64:27]
  assign _T_473 = _T_449 ? _T_472 : 13'h0; // @[Shift.scala 16:10]
  assign _T_474 = _T_473[12:12]; // @[convert.scala 23:34]
  assign decC_fraction = _T_473[11:0]; // @[convert.scala 24:34]
  assign _T_476 = _T_339 == 1'h0; // @[convert.scala 25:26]
  assign _T_478 = _T_339 ? _T_447 : _T_446; // @[convert.scala 25:42]
  assign _T_481 = ~ _T_474; // @[convert.scala 26:67]
  assign _T_482 = _T_337 ? _T_481 : _T_474; // @[convert.scala 26:51]
  assign _T_483 = {_T_476,_T_478,_T_482}; // @[Cat.scala 29:58]
  assign _T_485 = realC[14:0]; // @[convert.scala 29:56]
  assign _T_486 = _T_485 != 15'h0; // @[convert.scala 29:60]
  assign _T_487 = ~ _T_486; // @[convert.scala 29:41]
  assign decC_isNaR = _T_337 & _T_487; // @[convert.scala 29:39]
  assign _T_490 = _T_337 == 1'h0; // @[convert.scala 30:19]
  assign decC_isZero = _T_490 & _T_487; // @[convert.scala 30:41]
  assign decC_scale = $signed(_T_483); // @[convert.scala 32:24]
  assign _T_498 = decA_isNaR | decB_isNaR; // @[PositFMA.scala 58:30]
  assign outIsNaR = _T_498 | decC_isNaR; // @[PositFMA.scala 58:44]
  assign _T_499 = ~ _T_13; // @[PositFMA.scala 59:34]
  assign _T_500 = ~ decA_isZero; // @[PositFMA.scala 59:47]
  assign _T_501 = _T_499 & _T_500; // @[PositFMA.scala 59:45]
  assign _T_503 = {_T_13,_T_501,decA_fraction}; // @[Cat.scala 29:58]
  assign sigA = $signed(_T_503); // @[PositFMA.scala 59:76]
  assign _T_504 = ~ _T_175; // @[PositFMA.scala 60:34]
  assign _T_505 = ~ decB_isZero; // @[PositFMA.scala 60:47]
  assign _T_506 = _T_504 & _T_505; // @[PositFMA.scala 60:45]
  assign _T_508 = {_T_175,_T_506,decB_fraction}; // @[Cat.scala 29:58]
  assign sigB = $signed(_T_508); // @[PositFMA.scala 60:76]
  assign _T_509 = $signed(sigA) * $signed(sigB); // @[PositFMA.scala 61:25]
  assign sigP = $unsigned(_T_509); // @[PositFMA.scala 61:33]
  assign head2 = sigP[27:26]; // @[PositFMA.scala 62:28]
  assign _T_510 = head2[1]; // @[PositFMA.scala 63:31]
  assign _T_511 = ~ _T_510; // @[PositFMA.scala 63:25]
  assign _T_512 = head2[0]; // @[PositFMA.scala 63:42]
  assign addTwo = _T_511 & _T_512; // @[PositFMA.scala 63:35]
  assign _T_513 = sigP[27]; // @[PositFMA.scala 65:23]
  assign _T_514 = sigP[25]; // @[PositFMA.scala 65:49]
  assign addOne = _T_513 ^ _T_514; // @[PositFMA.scala 65:43]
  assign _T_515 = {addTwo,addOne}; // @[Cat.scala 29:58]
  assign expBias = {1'b0,$signed(_T_515)}; // @[PositFMA.scala 66:39]
  assign mulSign = sigP[27:27]; // @[PositFMA.scala 67:28]
  assign _T_516 = $signed(decA_scale) + $signed(decB_scale); // @[PositFMA.scala 69:30]
  assign _GEN_12 = {{4{expBias[2]}},expBias}; // @[PositFMA.scala 69:44]
  assign _T_518 = $signed(_T_516) + $signed(_GEN_12); // @[PositFMA.scala 69:44]
  assign mulScale = $signed(_T_518); // @[PositFMA.scala 69:44]
  assign _T_519 = sigP[25:0]; // @[PositFMA.scala 72:29]
  assign _T_520 = sigP[24:0]; // @[PositFMA.scala 73:29]
  assign _T_521 = {_T_520, 1'h0}; // @[PositFMA.scala 73:48]
  assign mulSigTmp = addOne ? _T_519 : _T_521; // @[PositFMA.scala 70:22]
  assign _T_523 = mulSigTmp[25:25]; // @[PositFMA.scala 77:39]
  assign _T_524 = _T_523 | addTwo; // @[PositFMA.scala 77:43]
  assign _T_525 = mulSigTmp[24:0]; // @[PositFMA.scala 78:39]
  assign mulSig = {mulSign,_T_524,_T_525}; // @[Cat.scala 29:58]
  assign _T_551 = ~ addSign_phase2; // @[PositFMA.scala 107:29]
  assign _T_552 = ~ addZero_phase2; // @[PositFMA.scala 107:47]
  assign _T_553 = _T_551 & _T_552; // @[PositFMA.scala 107:45]
  assign extAddSig = {addSign_phase2,_T_553,addFrac_phase2,13'h0}; // @[Cat.scala 29:58]
  assign _GEN_13 = {{1{addScale_phase2[5]}},addScale_phase2}; // @[PositFMA.scala 111:39]
  assign mulGreater = $signed(mulScale_phase2) > $signed(_GEN_13); // @[PositFMA.scala 111:39]
  assign greaterScale = mulGreater ? $signed(mulScale_phase2) : $signed({{1{addScale_phase2[5]}},addScale_phase2}); // @[PositFMA.scala 112:26]
  assign smallerScale = mulGreater ? $signed({{1{addScale_phase2[5]}},addScale_phase2}) : $signed(mulScale_phase2); // @[PositFMA.scala 113:26]
  assign _T_557 = $signed(greaterScale) - $signed(smallerScale); // @[PositFMA.scala 114:36]
  assign scaleDiff = $signed(_T_557); // @[PositFMA.scala 114:36]
  assign greaterSig = mulGreater ? mulSig_phase2 : extAddSig; // @[PositFMA.scala 115:26]
  assign smallerSigTmp = mulGreater ? extAddSig : mulSig_phase2; // @[PositFMA.scala 116:26]
  assign _T_558 = $unsigned(scaleDiff); // @[PositFMA.scala 117:69]
  assign _T_559 = _T_558 < 7'h1b; // @[Shift.scala 39:24]
  assign _T_560 = _T_558[4:0]; // @[Shift.scala 40:44]
  assign _T_561 = smallerSigTmp[26:16]; // @[Shift.scala 90:30]
  assign _T_562 = smallerSigTmp[15:0]; // @[Shift.scala 90:48]
  assign _T_563 = _T_562 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_14 = {{10'd0}, _T_563}; // @[Shift.scala 90:39]
  assign _T_564 = _T_561 | _GEN_14; // @[Shift.scala 90:39]
  assign _T_565 = _T_560[4]; // @[Shift.scala 12:21]
  assign _T_566 = smallerSigTmp[26]; // @[Shift.scala 12:21]
  assign _T_568 = _T_566 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_569 = {_T_568,_T_564}; // @[Cat.scala 29:58]
  assign _T_570 = _T_565 ? _T_569 : smallerSigTmp; // @[Shift.scala 91:22]
  assign _T_571 = _T_560[3:0]; // @[Shift.scala 92:77]
  assign _T_572 = _T_570[26:8]; // @[Shift.scala 90:30]
  assign _T_573 = _T_570[7:0]; // @[Shift.scala 90:48]
  assign _T_574 = _T_573 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_15 = {{18'd0}, _T_574}; // @[Shift.scala 90:39]
  assign _T_575 = _T_572 | _GEN_15; // @[Shift.scala 90:39]
  assign _T_576 = _T_571[3]; // @[Shift.scala 12:21]
  assign _T_577 = _T_570[26]; // @[Shift.scala 12:21]
  assign _T_579 = _T_577 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_580 = {_T_579,_T_575}; // @[Cat.scala 29:58]
  assign _T_581 = _T_576 ? _T_580 : _T_570; // @[Shift.scala 91:22]
  assign _T_582 = _T_571[2:0]; // @[Shift.scala 92:77]
  assign _T_583 = _T_581[26:4]; // @[Shift.scala 90:30]
  assign _T_584 = _T_581[3:0]; // @[Shift.scala 90:48]
  assign _T_585 = _T_584 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_16 = {{22'd0}, _T_585}; // @[Shift.scala 90:39]
  assign _T_586 = _T_583 | _GEN_16; // @[Shift.scala 90:39]
  assign _T_587 = _T_582[2]; // @[Shift.scala 12:21]
  assign _T_588 = _T_581[26]; // @[Shift.scala 12:21]
  assign _T_590 = _T_588 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_591 = {_T_590,_T_586}; // @[Cat.scala 29:58]
  assign _T_592 = _T_587 ? _T_591 : _T_581; // @[Shift.scala 91:22]
  assign _T_593 = _T_582[1:0]; // @[Shift.scala 92:77]
  assign _T_594 = _T_592[26:2]; // @[Shift.scala 90:30]
  assign _T_595 = _T_592[1:0]; // @[Shift.scala 90:48]
  assign _T_596 = _T_595 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_17 = {{24'd0}, _T_596}; // @[Shift.scala 90:39]
  assign _T_597 = _T_594 | _GEN_17; // @[Shift.scala 90:39]
  assign _T_598 = _T_593[1]; // @[Shift.scala 12:21]
  assign _T_599 = _T_592[26]; // @[Shift.scala 12:21]
  assign _T_601 = _T_599 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_602 = {_T_601,_T_597}; // @[Cat.scala 29:58]
  assign _T_603 = _T_598 ? _T_602 : _T_592; // @[Shift.scala 91:22]
  assign _T_604 = _T_593[0:0]; // @[Shift.scala 92:77]
  assign _T_605 = _T_603[26:1]; // @[Shift.scala 90:30]
  assign _T_606 = _T_603[0:0]; // @[Shift.scala 90:48]
  assign _GEN_18 = {{25'd0}, _T_606}; // @[Shift.scala 90:39]
  assign _T_608 = _T_605 | _GEN_18; // @[Shift.scala 90:39]
  assign _T_610 = _T_603[26]; // @[Shift.scala 12:21]
  assign _T_611 = {_T_610,_T_608}; // @[Cat.scala 29:58]
  assign _T_612 = _T_604 ? _T_611 : _T_603; // @[Shift.scala 91:22]
  assign _T_615 = _T_566 ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_559 ? _T_612 : _T_615; // @[Shift.scala 39:10]
  assign rawSumSig = greaterSig + smallerSig; // @[PositFMA.scala 118:34]
  assign _T_616 = mulSig_phase2[26:26]; // @[PositFMA.scala 119:42]
  assign _T_617 = _T_616 ^ addSign_phase2; // @[PositFMA.scala 119:46]
  assign _T_618 = rawSumSig[27:27]; // @[PositFMA.scala 119:79]
  assign sumSign = _T_617 ^ _T_618; // @[PositFMA.scala 119:63]
  assign _T_620 = greaterSig + smallerSig; // @[PositFMA.scala 120:50]
  assign signSumSig = {sumSign,_T_620}; // @[Cat.scala 29:58]
  assign _T_621 = signSumSig[27:1]; // @[PositFMA.scala 124:33]
  assign _T_622 = signSumSig[26:0]; // @[PositFMA.scala 124:68]
  assign sumXor = _T_621 ^ _T_622; // @[PositFMA.scala 124:51]
  assign _T_623 = sumXor[26:11]; // @[LZD.scala 43:32]
  assign _T_624 = _T_623[15:8]; // @[LZD.scala 43:32]
  assign _T_625 = _T_624[7:4]; // @[LZD.scala 43:32]
  assign _T_626 = _T_625[3:2]; // @[LZD.scala 43:32]
  assign _T_627 = _T_626 != 2'h0; // @[LZD.scala 39:14]
  assign _T_628 = _T_626[1]; // @[LZD.scala 39:21]
  assign _T_629 = _T_626[0]; // @[LZD.scala 39:30]
  assign _T_630 = ~ _T_629; // @[LZD.scala 39:27]
  assign _T_631 = _T_628 | _T_630; // @[LZD.scala 39:25]
  assign _T_632 = {_T_627,_T_631}; // @[Cat.scala 29:58]
  assign _T_633 = _T_625[1:0]; // @[LZD.scala 44:32]
  assign _T_634 = _T_633 != 2'h0; // @[LZD.scala 39:14]
  assign _T_635 = _T_633[1]; // @[LZD.scala 39:21]
  assign _T_636 = _T_633[0]; // @[LZD.scala 39:30]
  assign _T_637 = ~ _T_636; // @[LZD.scala 39:27]
  assign _T_638 = _T_635 | _T_637; // @[LZD.scala 39:25]
  assign _T_639 = {_T_634,_T_638}; // @[Cat.scala 29:58]
  assign _T_640 = _T_632[1]; // @[Shift.scala 12:21]
  assign _T_641 = _T_639[1]; // @[Shift.scala 12:21]
  assign _T_642 = _T_640 | _T_641; // @[LZD.scala 49:16]
  assign _T_643 = ~ _T_641; // @[LZD.scala 49:27]
  assign _T_644 = _T_640 | _T_643; // @[LZD.scala 49:25]
  assign _T_645 = _T_632[0:0]; // @[LZD.scala 49:47]
  assign _T_646 = _T_639[0:0]; // @[LZD.scala 49:59]
  assign _T_647 = _T_640 ? _T_645 : _T_646; // @[LZD.scala 49:35]
  assign _T_649 = {_T_642,_T_644,_T_647}; // @[Cat.scala 29:58]
  assign _T_650 = _T_624[3:0]; // @[LZD.scala 44:32]
  assign _T_651 = _T_650[3:2]; // @[LZD.scala 43:32]
  assign _T_652 = _T_651 != 2'h0; // @[LZD.scala 39:14]
  assign _T_653 = _T_651[1]; // @[LZD.scala 39:21]
  assign _T_654 = _T_651[0]; // @[LZD.scala 39:30]
  assign _T_655 = ~ _T_654; // @[LZD.scala 39:27]
  assign _T_656 = _T_653 | _T_655; // @[LZD.scala 39:25]
  assign _T_657 = {_T_652,_T_656}; // @[Cat.scala 29:58]
  assign _T_658 = _T_650[1:0]; // @[LZD.scala 44:32]
  assign _T_659 = _T_658 != 2'h0; // @[LZD.scala 39:14]
  assign _T_660 = _T_658[1]; // @[LZD.scala 39:21]
  assign _T_661 = _T_658[0]; // @[LZD.scala 39:30]
  assign _T_662 = ~ _T_661; // @[LZD.scala 39:27]
  assign _T_663 = _T_660 | _T_662; // @[LZD.scala 39:25]
  assign _T_664 = {_T_659,_T_663}; // @[Cat.scala 29:58]
  assign _T_665 = _T_657[1]; // @[Shift.scala 12:21]
  assign _T_666 = _T_664[1]; // @[Shift.scala 12:21]
  assign _T_667 = _T_665 | _T_666; // @[LZD.scala 49:16]
  assign _T_668 = ~ _T_666; // @[LZD.scala 49:27]
  assign _T_669 = _T_665 | _T_668; // @[LZD.scala 49:25]
  assign _T_670 = _T_657[0:0]; // @[LZD.scala 49:47]
  assign _T_671 = _T_664[0:0]; // @[LZD.scala 49:59]
  assign _T_672 = _T_665 ? _T_670 : _T_671; // @[LZD.scala 49:35]
  assign _T_674 = {_T_667,_T_669,_T_672}; // @[Cat.scala 29:58]
  assign _T_675 = _T_649[2]; // @[Shift.scala 12:21]
  assign _T_676 = _T_674[2]; // @[Shift.scala 12:21]
  assign _T_677 = _T_675 | _T_676; // @[LZD.scala 49:16]
  assign _T_678 = ~ _T_676; // @[LZD.scala 49:27]
  assign _T_679 = _T_675 | _T_678; // @[LZD.scala 49:25]
  assign _T_680 = _T_649[1:0]; // @[LZD.scala 49:47]
  assign _T_681 = _T_674[1:0]; // @[LZD.scala 49:59]
  assign _T_682 = _T_675 ? _T_680 : _T_681; // @[LZD.scala 49:35]
  assign _T_684 = {_T_677,_T_679,_T_682}; // @[Cat.scala 29:58]
  assign _T_685 = _T_623[7:0]; // @[LZD.scala 44:32]
  assign _T_686 = _T_685[7:4]; // @[LZD.scala 43:32]
  assign _T_687 = _T_686[3:2]; // @[LZD.scala 43:32]
  assign _T_688 = _T_687 != 2'h0; // @[LZD.scala 39:14]
  assign _T_689 = _T_687[1]; // @[LZD.scala 39:21]
  assign _T_690 = _T_687[0]; // @[LZD.scala 39:30]
  assign _T_691 = ~ _T_690; // @[LZD.scala 39:27]
  assign _T_692 = _T_689 | _T_691; // @[LZD.scala 39:25]
  assign _T_693 = {_T_688,_T_692}; // @[Cat.scala 29:58]
  assign _T_694 = _T_686[1:0]; // @[LZD.scala 44:32]
  assign _T_695 = _T_694 != 2'h0; // @[LZD.scala 39:14]
  assign _T_696 = _T_694[1]; // @[LZD.scala 39:21]
  assign _T_697 = _T_694[0]; // @[LZD.scala 39:30]
  assign _T_698 = ~ _T_697; // @[LZD.scala 39:27]
  assign _T_699 = _T_696 | _T_698; // @[LZD.scala 39:25]
  assign _T_700 = {_T_695,_T_699}; // @[Cat.scala 29:58]
  assign _T_701 = _T_693[1]; // @[Shift.scala 12:21]
  assign _T_702 = _T_700[1]; // @[Shift.scala 12:21]
  assign _T_703 = _T_701 | _T_702; // @[LZD.scala 49:16]
  assign _T_704 = ~ _T_702; // @[LZD.scala 49:27]
  assign _T_705 = _T_701 | _T_704; // @[LZD.scala 49:25]
  assign _T_706 = _T_693[0:0]; // @[LZD.scala 49:47]
  assign _T_707 = _T_700[0:0]; // @[LZD.scala 49:59]
  assign _T_708 = _T_701 ? _T_706 : _T_707; // @[LZD.scala 49:35]
  assign _T_710 = {_T_703,_T_705,_T_708}; // @[Cat.scala 29:58]
  assign _T_711 = _T_685[3:0]; // @[LZD.scala 44:32]
  assign _T_712 = _T_711[3:2]; // @[LZD.scala 43:32]
  assign _T_713 = _T_712 != 2'h0; // @[LZD.scala 39:14]
  assign _T_714 = _T_712[1]; // @[LZD.scala 39:21]
  assign _T_715 = _T_712[0]; // @[LZD.scala 39:30]
  assign _T_716 = ~ _T_715; // @[LZD.scala 39:27]
  assign _T_717 = _T_714 | _T_716; // @[LZD.scala 39:25]
  assign _T_718 = {_T_713,_T_717}; // @[Cat.scala 29:58]
  assign _T_719 = _T_711[1:0]; // @[LZD.scala 44:32]
  assign _T_720 = _T_719 != 2'h0; // @[LZD.scala 39:14]
  assign _T_721 = _T_719[1]; // @[LZD.scala 39:21]
  assign _T_722 = _T_719[0]; // @[LZD.scala 39:30]
  assign _T_723 = ~ _T_722; // @[LZD.scala 39:27]
  assign _T_724 = _T_721 | _T_723; // @[LZD.scala 39:25]
  assign _T_725 = {_T_720,_T_724}; // @[Cat.scala 29:58]
  assign _T_726 = _T_718[1]; // @[Shift.scala 12:21]
  assign _T_727 = _T_725[1]; // @[Shift.scala 12:21]
  assign _T_728 = _T_726 | _T_727; // @[LZD.scala 49:16]
  assign _T_729 = ~ _T_727; // @[LZD.scala 49:27]
  assign _T_730 = _T_726 | _T_729; // @[LZD.scala 49:25]
  assign _T_731 = _T_718[0:0]; // @[LZD.scala 49:47]
  assign _T_732 = _T_725[0:0]; // @[LZD.scala 49:59]
  assign _T_733 = _T_726 ? _T_731 : _T_732; // @[LZD.scala 49:35]
  assign _T_735 = {_T_728,_T_730,_T_733}; // @[Cat.scala 29:58]
  assign _T_736 = _T_710[2]; // @[Shift.scala 12:21]
  assign _T_737 = _T_735[2]; // @[Shift.scala 12:21]
  assign _T_738 = _T_736 | _T_737; // @[LZD.scala 49:16]
  assign _T_739 = ~ _T_737; // @[LZD.scala 49:27]
  assign _T_740 = _T_736 | _T_739; // @[LZD.scala 49:25]
  assign _T_741 = _T_710[1:0]; // @[LZD.scala 49:47]
  assign _T_742 = _T_735[1:0]; // @[LZD.scala 49:59]
  assign _T_743 = _T_736 ? _T_741 : _T_742; // @[LZD.scala 49:35]
  assign _T_745 = {_T_738,_T_740,_T_743}; // @[Cat.scala 29:58]
  assign _T_746 = _T_684[3]; // @[Shift.scala 12:21]
  assign _T_747 = _T_745[3]; // @[Shift.scala 12:21]
  assign _T_748 = _T_746 | _T_747; // @[LZD.scala 49:16]
  assign _T_749 = ~ _T_747; // @[LZD.scala 49:27]
  assign _T_750 = _T_746 | _T_749; // @[LZD.scala 49:25]
  assign _T_751 = _T_684[2:0]; // @[LZD.scala 49:47]
  assign _T_752 = _T_745[2:0]; // @[LZD.scala 49:59]
  assign _T_753 = _T_746 ? _T_751 : _T_752; // @[LZD.scala 49:35]
  assign _T_755 = {_T_748,_T_750,_T_753}; // @[Cat.scala 29:58]
  assign _T_756 = sumXor[10:0]; // @[LZD.scala 44:32]
  assign _T_757 = _T_756[10:3]; // @[LZD.scala 43:32]
  assign _T_758 = _T_757[7:4]; // @[LZD.scala 43:32]
  assign _T_759 = _T_758[3:2]; // @[LZD.scala 43:32]
  assign _T_760 = _T_759 != 2'h0; // @[LZD.scala 39:14]
  assign _T_761 = _T_759[1]; // @[LZD.scala 39:21]
  assign _T_762 = _T_759[0]; // @[LZD.scala 39:30]
  assign _T_763 = ~ _T_762; // @[LZD.scala 39:27]
  assign _T_764 = _T_761 | _T_763; // @[LZD.scala 39:25]
  assign _T_765 = {_T_760,_T_764}; // @[Cat.scala 29:58]
  assign _T_766 = _T_758[1:0]; // @[LZD.scala 44:32]
  assign _T_767 = _T_766 != 2'h0; // @[LZD.scala 39:14]
  assign _T_768 = _T_766[1]; // @[LZD.scala 39:21]
  assign _T_769 = _T_766[0]; // @[LZD.scala 39:30]
  assign _T_770 = ~ _T_769; // @[LZD.scala 39:27]
  assign _T_771 = _T_768 | _T_770; // @[LZD.scala 39:25]
  assign _T_772 = {_T_767,_T_771}; // @[Cat.scala 29:58]
  assign _T_773 = _T_765[1]; // @[Shift.scala 12:21]
  assign _T_774 = _T_772[1]; // @[Shift.scala 12:21]
  assign _T_775 = _T_773 | _T_774; // @[LZD.scala 49:16]
  assign _T_776 = ~ _T_774; // @[LZD.scala 49:27]
  assign _T_777 = _T_773 | _T_776; // @[LZD.scala 49:25]
  assign _T_778 = _T_765[0:0]; // @[LZD.scala 49:47]
  assign _T_779 = _T_772[0:0]; // @[LZD.scala 49:59]
  assign _T_780 = _T_773 ? _T_778 : _T_779; // @[LZD.scala 49:35]
  assign _T_782 = {_T_775,_T_777,_T_780}; // @[Cat.scala 29:58]
  assign _T_783 = _T_757[3:0]; // @[LZD.scala 44:32]
  assign _T_784 = _T_783[3:2]; // @[LZD.scala 43:32]
  assign _T_785 = _T_784 != 2'h0; // @[LZD.scala 39:14]
  assign _T_786 = _T_784[1]; // @[LZD.scala 39:21]
  assign _T_787 = _T_784[0]; // @[LZD.scala 39:30]
  assign _T_788 = ~ _T_787; // @[LZD.scala 39:27]
  assign _T_789 = _T_786 | _T_788; // @[LZD.scala 39:25]
  assign _T_790 = {_T_785,_T_789}; // @[Cat.scala 29:58]
  assign _T_791 = _T_783[1:0]; // @[LZD.scala 44:32]
  assign _T_792 = _T_791 != 2'h0; // @[LZD.scala 39:14]
  assign _T_793 = _T_791[1]; // @[LZD.scala 39:21]
  assign _T_794 = _T_791[0]; // @[LZD.scala 39:30]
  assign _T_795 = ~ _T_794; // @[LZD.scala 39:27]
  assign _T_796 = _T_793 | _T_795; // @[LZD.scala 39:25]
  assign _T_797 = {_T_792,_T_796}; // @[Cat.scala 29:58]
  assign _T_798 = _T_790[1]; // @[Shift.scala 12:21]
  assign _T_799 = _T_797[1]; // @[Shift.scala 12:21]
  assign _T_800 = _T_798 | _T_799; // @[LZD.scala 49:16]
  assign _T_801 = ~ _T_799; // @[LZD.scala 49:27]
  assign _T_802 = _T_798 | _T_801; // @[LZD.scala 49:25]
  assign _T_803 = _T_790[0:0]; // @[LZD.scala 49:47]
  assign _T_804 = _T_797[0:0]; // @[LZD.scala 49:59]
  assign _T_805 = _T_798 ? _T_803 : _T_804; // @[LZD.scala 49:35]
  assign _T_807 = {_T_800,_T_802,_T_805}; // @[Cat.scala 29:58]
  assign _T_808 = _T_782[2]; // @[Shift.scala 12:21]
  assign _T_809 = _T_807[2]; // @[Shift.scala 12:21]
  assign _T_810 = _T_808 | _T_809; // @[LZD.scala 49:16]
  assign _T_811 = ~ _T_809; // @[LZD.scala 49:27]
  assign _T_812 = _T_808 | _T_811; // @[LZD.scala 49:25]
  assign _T_813 = _T_782[1:0]; // @[LZD.scala 49:47]
  assign _T_814 = _T_807[1:0]; // @[LZD.scala 49:59]
  assign _T_815 = _T_808 ? _T_813 : _T_814; // @[LZD.scala 49:35]
  assign _T_817 = {_T_810,_T_812,_T_815}; // @[Cat.scala 29:58]
  assign _T_818 = _T_756[2:0]; // @[LZD.scala 44:32]
  assign _T_819 = _T_818[2:1]; // @[LZD.scala 43:32]
  assign _T_820 = _T_819 != 2'h0; // @[LZD.scala 39:14]
  assign _T_821 = _T_819[1]; // @[LZD.scala 39:21]
  assign _T_822 = _T_819[0]; // @[LZD.scala 39:30]
  assign _T_823 = ~ _T_822; // @[LZD.scala 39:27]
  assign _T_824 = _T_821 | _T_823; // @[LZD.scala 39:25]
  assign _T_825 = {_T_820,_T_824}; // @[Cat.scala 29:58]
  assign _T_826 = _T_818[0:0]; // @[LZD.scala 44:32]
  assign _T_828 = _T_825[1]; // @[Shift.scala 12:21]
  assign _T_830 = _T_825[0:0]; // @[LZD.scala 55:32]
  assign _T_831 = _T_828 ? _T_830 : _T_826; // @[LZD.scala 55:20]
  assign _T_833 = _T_817[3]; // @[Shift.scala 12:21]
  assign _T_835 = {1'h1,_T_828,_T_831}; // @[Cat.scala 29:58]
  assign _T_836 = _T_817[2:0]; // @[LZD.scala 55:32]
  assign _T_837 = _T_833 ? _T_836 : _T_835; // @[LZD.scala 55:20]
  assign _T_838 = {_T_833,_T_837}; // @[Cat.scala 29:58]
  assign _T_839 = _T_755[4]; // @[Shift.scala 12:21]
  assign _T_841 = _T_755[3:0]; // @[LZD.scala 55:32]
  assign _T_842 = _T_839 ? _T_841 : _T_838; // @[LZD.scala 55:20]
  assign sumLZD = {_T_839,_T_842}; // @[Cat.scala 29:58]
  assign shiftValue = ~ sumLZD; // @[PositFMA.scala 126:24]
  assign _T_843 = signSumSig[25:0]; // @[PositFMA.scala 127:38]
  assign _T_844 = shiftValue < 5'h1a; // @[Shift.scala 16:24]
  assign _T_846 = shiftValue[4]; // @[Shift.scala 12:21]
  assign _T_847 = _T_843[9:0]; // @[Shift.scala 64:52]
  assign _T_849 = {_T_847,16'h0}; // @[Cat.scala 29:58]
  assign _T_850 = _T_846 ? _T_849 : _T_843; // @[Shift.scala 64:27]
  assign _T_851 = shiftValue[3:0]; // @[Shift.scala 66:70]
  assign _T_852 = _T_851[3]; // @[Shift.scala 12:21]
  assign _T_853 = _T_850[17:0]; // @[Shift.scala 64:52]
  assign _T_855 = {_T_853,8'h0}; // @[Cat.scala 29:58]
  assign _T_856 = _T_852 ? _T_855 : _T_850; // @[Shift.scala 64:27]
  assign _T_857 = _T_851[2:0]; // @[Shift.scala 66:70]
  assign _T_858 = _T_857[2]; // @[Shift.scala 12:21]
  assign _T_859 = _T_856[21:0]; // @[Shift.scala 64:52]
  assign _T_861 = {_T_859,4'h0}; // @[Cat.scala 29:58]
  assign _T_862 = _T_858 ? _T_861 : _T_856; // @[Shift.scala 64:27]
  assign _T_863 = _T_857[1:0]; // @[Shift.scala 66:70]
  assign _T_864 = _T_863[1]; // @[Shift.scala 12:21]
  assign _T_865 = _T_862[23:0]; // @[Shift.scala 64:52]
  assign _T_867 = {_T_865,2'h0}; // @[Cat.scala 29:58]
  assign _T_868 = _T_864 ? _T_867 : _T_862; // @[Shift.scala 64:27]
  assign _T_869 = _T_863[0:0]; // @[Shift.scala 66:70]
  assign _T_871 = _T_868[24:0]; // @[Shift.scala 64:52]
  assign _T_872 = {_T_871,1'h0}; // @[Cat.scala 29:58]
  assign _T_873 = _T_869 ? _T_872 : _T_868; // @[Shift.scala 64:27]
  assign normalFracTmp = _T_844 ? _T_873 : 26'h0; // @[Shift.scala 16:10]
  assign _T_875 = $signed(greaterScale) + $signed(7'sh2); // @[PositFMA.scala 130:36]
  assign _T_876 = $signed(_T_875); // @[PositFMA.scala 130:36]
  assign _T_877 = {1'h1,_T_839,_T_842}; // @[Cat.scala 29:58]
  assign _T_878 = $signed(_T_877); // @[PositFMA.scala 130:61]
  assign _GEN_19 = {{1{_T_878[5]}},_T_878}; // @[PositFMA.scala 130:42]
  assign _T_880 = $signed(_T_876) + $signed(_GEN_19); // @[PositFMA.scala 130:42]
  assign sumScale = $signed(_T_880); // @[PositFMA.scala 130:42]
  assign sumFrac = normalFracTmp[25:14]; // @[PositFMA.scala 131:41]
  assign grsTmp = normalFracTmp[13:0]; // @[PositFMA.scala 134:41]
  assign _T_881 = grsTmp[13:12]; // @[PositFMA.scala 137:40]
  assign _T_882 = grsTmp[11:0]; // @[PositFMA.scala 137:56]
  assign _T_883 = _T_882 != 12'h0; // @[PositFMA.scala 137:60]
  assign underflow = $signed(sumScale) < $signed(-7'sh1d); // @[PositFMA.scala 144:32]
  assign overflow = $signed(sumScale) > $signed(7'sh1c); // @[PositFMA.scala 145:32]
  assign _T_884 = signSumSig != 28'h0; // @[PositFMA.scala 154:32]
  assign decF_isZero = ~ _T_884; // @[PositFMA.scala 154:20]
  assign _T_886 = underflow ? $signed(-7'sh1d) : $signed(sumScale); // @[Mux.scala 87:16]
  assign _T_887 = overflow ? $signed(7'sh1c) : $signed(_T_886); // @[Mux.scala 87:16]
  assign _GEN_20 = _T_887[5:0]; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  assign decF_scale = $signed(_GEN_20); // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  assign _T_888 = decF_scale[0]; // @[convert.scala 46:61]
  assign _T_889 = ~ _T_888; // @[convert.scala 46:52]
  assign _T_891 = sumSign ? _T_889 : _T_888; // @[convert.scala 46:42]
  assign _T_892 = decF_scale[5:1]; // @[convert.scala 48:34]
  assign _T_893 = _T_892[4:4]; // @[convert.scala 49:36]
  assign _T_895 = ~ _T_892; // @[convert.scala 50:36]
  assign _T_896 = $signed(_T_895); // @[convert.scala 50:36]
  assign _T_897 = _T_893 ? $signed(_T_896) : $signed(_T_892); // @[convert.scala 50:28]
  assign _T_898 = _T_893 ^ sumSign; // @[convert.scala 51:31]
  assign _T_899 = ~ _T_898; // @[convert.scala 52:43]
  assign _T_903 = {_T_899,_T_898,_T_891,sumFrac,_T_881,_T_883}; // @[Cat.scala 29:58]
  assign _T_904 = $unsigned(_T_897); // @[Shift.scala 39:17]
  assign _T_905 = _T_904 < 5'h12; // @[Shift.scala 39:24]
  assign _T_907 = _T_903[17:16]; // @[Shift.scala 90:30]
  assign _T_908 = _T_903[15:0]; // @[Shift.scala 90:48]
  assign _T_909 = _T_908 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_21 = {{1'd0}, _T_909}; // @[Shift.scala 90:39]
  assign _T_910 = _T_907 | _GEN_21; // @[Shift.scala 90:39]
  assign _T_911 = _T_904[4]; // @[Shift.scala 12:21]
  assign _T_912 = _T_903[17]; // @[Shift.scala 12:21]
  assign _T_914 = _T_912 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_915 = {_T_914,_T_910}; // @[Cat.scala 29:58]
  assign _T_916 = _T_911 ? _T_915 : _T_903; // @[Shift.scala 91:22]
  assign _T_917 = _T_904[3:0]; // @[Shift.scala 92:77]
  assign _T_918 = _T_916[17:8]; // @[Shift.scala 90:30]
  assign _T_919 = _T_916[7:0]; // @[Shift.scala 90:48]
  assign _T_920 = _T_919 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_22 = {{9'd0}, _T_920}; // @[Shift.scala 90:39]
  assign _T_921 = _T_918 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_922 = _T_917[3]; // @[Shift.scala 12:21]
  assign _T_923 = _T_916[17]; // @[Shift.scala 12:21]
  assign _T_925 = _T_923 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_926 = {_T_925,_T_921}; // @[Cat.scala 29:58]
  assign _T_927 = _T_922 ? _T_926 : _T_916; // @[Shift.scala 91:22]
  assign _T_928 = _T_917[2:0]; // @[Shift.scala 92:77]
  assign _T_929 = _T_927[17:4]; // @[Shift.scala 90:30]
  assign _T_930 = _T_927[3:0]; // @[Shift.scala 90:48]
  assign _T_931 = _T_930 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_23 = {{13'd0}, _T_931}; // @[Shift.scala 90:39]
  assign _T_932 = _T_929 | _GEN_23; // @[Shift.scala 90:39]
  assign _T_933 = _T_928[2]; // @[Shift.scala 12:21]
  assign _T_934 = _T_927[17]; // @[Shift.scala 12:21]
  assign _T_936 = _T_934 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_937 = {_T_936,_T_932}; // @[Cat.scala 29:58]
  assign _T_938 = _T_933 ? _T_937 : _T_927; // @[Shift.scala 91:22]
  assign _T_939 = _T_928[1:0]; // @[Shift.scala 92:77]
  assign _T_940 = _T_938[17:2]; // @[Shift.scala 90:30]
  assign _T_941 = _T_938[1:0]; // @[Shift.scala 90:48]
  assign _T_942 = _T_941 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_24 = {{15'd0}, _T_942}; // @[Shift.scala 90:39]
  assign _T_943 = _T_940 | _GEN_24; // @[Shift.scala 90:39]
  assign _T_944 = _T_939[1]; // @[Shift.scala 12:21]
  assign _T_945 = _T_938[17]; // @[Shift.scala 12:21]
  assign _T_947 = _T_945 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_948 = {_T_947,_T_943}; // @[Cat.scala 29:58]
  assign _T_949 = _T_944 ? _T_948 : _T_938; // @[Shift.scala 91:22]
  assign _T_950 = _T_939[0:0]; // @[Shift.scala 92:77]
  assign _T_951 = _T_949[17:1]; // @[Shift.scala 90:30]
  assign _T_952 = _T_949[0:0]; // @[Shift.scala 90:48]
  assign _GEN_25 = {{16'd0}, _T_952}; // @[Shift.scala 90:39]
  assign _T_954 = _T_951 | _GEN_25; // @[Shift.scala 90:39]
  assign _T_956 = _T_949[17]; // @[Shift.scala 12:21]
  assign _T_957 = {_T_956,_T_954}; // @[Cat.scala 29:58]
  assign _T_958 = _T_950 ? _T_957 : _T_949; // @[Shift.scala 91:22]
  assign _T_961 = _T_912 ? 18'h3ffff : 18'h0; // @[Bitwise.scala 71:12]
  assign _T_962 = _T_905 ? _T_958 : _T_961; // @[Shift.scala 39:10]
  assign _T_963 = _T_962[3]; // @[convert.scala 55:31]
  assign _T_964 = _T_962[2]; // @[convert.scala 56:31]
  assign _T_965 = _T_962[1]; // @[convert.scala 57:31]
  assign _T_966 = _T_962[0]; // @[convert.scala 58:31]
  assign _T_967 = _T_962[17:3]; // @[convert.scala 59:69]
  assign _T_968 = _T_967 != 15'h0; // @[convert.scala 59:81]
  assign _T_969 = ~ _T_968; // @[convert.scala 59:50]
  assign _T_971 = _T_967 == 15'h7fff; // @[convert.scala 60:81]
  assign _T_972 = _T_963 | _T_965; // @[convert.scala 61:44]
  assign _T_973 = _T_972 | _T_966; // @[convert.scala 61:52]
  assign _T_974 = _T_964 & _T_973; // @[convert.scala 61:36]
  assign _T_975 = ~ _T_971; // @[convert.scala 62:63]
  assign _T_976 = _T_975 & _T_974; // @[convert.scala 62:103]
  assign _T_977 = _T_969 | _T_976; // @[convert.scala 62:60]
  assign _GEN_26 = {{14'd0}, _T_977}; // @[convert.scala 63:56]
  assign _T_980 = _T_967 + _GEN_26; // @[convert.scala 63:56]
  assign _T_981 = {sumSign,_T_980}; // @[Cat.scala 29:58]
  assign io_F = _T_989; // @[PositFMA.scala 174:15]
  assign io_outValid = _T_985; // @[PositFMA.scala 173:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  outIsNaR_phase2 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mulSig_phase2 = _RAND_1[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  addFrac_phase2 = _RAND_2[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mulScale_phase2 = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addScale_phase2 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addSign_phase2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addZero_phase2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  inValid_phase2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_985 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_989 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (io_inValid) begin
      outIsNaR_phase2 <= outIsNaR;
    end
    if (io_inValid) begin
      mulSig_phase2 <= mulSig;
    end
    if (io_inValid) begin
      addFrac_phase2 <= decC_fraction;
    end
    if (io_inValid) begin
      mulScale_phase2 <= mulScale;
    end
    if (io_inValid) begin
      addScale_phase2 <= decC_scale;
    end
    if (io_inValid) begin
      addSign_phase2 <= _T_337;
    end
    if (io_inValid) begin
      addZero_phase2 <= decC_isZero;
    end
    if (reset) begin
      inValid_phase2 <= 1'h0;
    end else begin
      inValid_phase2 <= io_inValid;
    end
    if (reset) begin
      _T_985 <= 1'h0;
    end else begin
      _T_985 <= inValid_phase2;
    end
    if (inValid_phase2) begin
      if (outIsNaR_phase2) begin
        _T_989 <= 16'h8000;
      end else begin
        if (decF_isZero) begin
          _T_989 <= 16'h0;
        end else begin
          _T_989 <= _T_981;
        end
      end
    end
  end
endmodule
