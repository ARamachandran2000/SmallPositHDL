module PositFMA32_1(
  input         clock,
  input         reset,
  input         io_inValid,
  input  [1:0]  io_fmaOp,
  input  [31:0] io_A,
  input  [31:0] io_B,
  input  [31:0] io_C,
  output [31:0] io_F,
  output        io_outValid
);
  wire  _T; // @[PositFMA.scala 47:36]
  wire [31:0] _T_2; // @[Bitwise.scala 71:12]
  wire [31:0] _T_3; // @[PositFMA.scala 47:41]
  wire [31:0] _GEN_10; // @[PositFMA.scala 47:49]
  wire [31:0] realA; // @[PositFMA.scala 47:49]
  wire  _T_6; // @[PositFMA.scala 48:36]
  wire [31:0] _T_8; // @[Bitwise.scala 71:12]
  wire [31:0] _T_9; // @[PositFMA.scala 48:41]
  wire [31:0] _GEN_11; // @[PositFMA.scala 48:49]
  wire [31:0] realC; // @[PositFMA.scala 48:49]
  wire  _T_13; // @[convert.scala 18:24]
  wire  _T_14; // @[convert.scala 18:40]
  wire  _T_15; // @[convert.scala 18:36]
  wire [29:0] _T_16; // @[convert.scala 19:24]
  wire [29:0] _T_17; // @[convert.scala 19:43]
  wire [29:0] _T_18; // @[convert.scala 19:39]
  wire [15:0] _T_19; // @[LZD.scala 43:32]
  wire [7:0] _T_20; // @[LZD.scala 43:32]
  wire [3:0] _T_21; // @[LZD.scala 43:32]
  wire [1:0] _T_22; // @[LZD.scala 43:32]
  wire  _T_23; // @[LZD.scala 39:14]
  wire  _T_24; // @[LZD.scala 39:21]
  wire  _T_25; // @[LZD.scala 39:30]
  wire  _T_26; // @[LZD.scala 39:27]
  wire  _T_27; // @[LZD.scala 39:25]
  wire [1:0] _T_28; // @[Cat.scala 29:58]
  wire [1:0] _T_29; // @[LZD.scala 44:32]
  wire  _T_30; // @[LZD.scala 39:14]
  wire  _T_31; // @[LZD.scala 39:21]
  wire  _T_32; // @[LZD.scala 39:30]
  wire  _T_33; // @[LZD.scala 39:27]
  wire  _T_34; // @[LZD.scala 39:25]
  wire [1:0] _T_35; // @[Cat.scala 29:58]
  wire  _T_36; // @[Shift.scala 12:21]
  wire  _T_37; // @[Shift.scala 12:21]
  wire  _T_38; // @[LZD.scala 49:16]
  wire  _T_39; // @[LZD.scala 49:27]
  wire  _T_40; // @[LZD.scala 49:25]
  wire  _T_41; // @[LZD.scala 49:47]
  wire  _T_42; // @[LZD.scala 49:59]
  wire  _T_43; // @[LZD.scala 49:35]
  wire [2:0] _T_45; // @[Cat.scala 29:58]
  wire [3:0] _T_46; // @[LZD.scala 44:32]
  wire [1:0] _T_47; // @[LZD.scala 43:32]
  wire  _T_48; // @[LZD.scala 39:14]
  wire  _T_49; // @[LZD.scala 39:21]
  wire  _T_50; // @[LZD.scala 39:30]
  wire  _T_51; // @[LZD.scala 39:27]
  wire  _T_52; // @[LZD.scala 39:25]
  wire [1:0] _T_53; // @[Cat.scala 29:58]
  wire [1:0] _T_54; // @[LZD.scala 44:32]
  wire  _T_55; // @[LZD.scala 39:14]
  wire  _T_56; // @[LZD.scala 39:21]
  wire  _T_57; // @[LZD.scala 39:30]
  wire  _T_58; // @[LZD.scala 39:27]
  wire  _T_59; // @[LZD.scala 39:25]
  wire [1:0] _T_60; // @[Cat.scala 29:58]
  wire  _T_61; // @[Shift.scala 12:21]
  wire  _T_62; // @[Shift.scala 12:21]
  wire  _T_63; // @[LZD.scala 49:16]
  wire  _T_64; // @[LZD.scala 49:27]
  wire  _T_65; // @[LZD.scala 49:25]
  wire  _T_66; // @[LZD.scala 49:47]
  wire  _T_67; // @[LZD.scala 49:59]
  wire  _T_68; // @[LZD.scala 49:35]
  wire [2:0] _T_70; // @[Cat.scala 29:58]
  wire  _T_71; // @[Shift.scala 12:21]
  wire  _T_72; // @[Shift.scala 12:21]
  wire  _T_73; // @[LZD.scala 49:16]
  wire  _T_74; // @[LZD.scala 49:27]
  wire  _T_75; // @[LZD.scala 49:25]
  wire [1:0] _T_76; // @[LZD.scala 49:47]
  wire [1:0] _T_77; // @[LZD.scala 49:59]
  wire [1:0] _T_78; // @[LZD.scala 49:35]
  wire [3:0] _T_80; // @[Cat.scala 29:58]
  wire [7:0] _T_81; // @[LZD.scala 44:32]
  wire [3:0] _T_82; // @[LZD.scala 43:32]
  wire [1:0] _T_83; // @[LZD.scala 43:32]
  wire  _T_84; // @[LZD.scala 39:14]
  wire  _T_85; // @[LZD.scala 39:21]
  wire  _T_86; // @[LZD.scala 39:30]
  wire  _T_87; // @[LZD.scala 39:27]
  wire  _T_88; // @[LZD.scala 39:25]
  wire [1:0] _T_89; // @[Cat.scala 29:58]
  wire [1:0] _T_90; // @[LZD.scala 44:32]
  wire  _T_91; // @[LZD.scala 39:14]
  wire  _T_92; // @[LZD.scala 39:21]
  wire  _T_93; // @[LZD.scala 39:30]
  wire  _T_94; // @[LZD.scala 39:27]
  wire  _T_95; // @[LZD.scala 39:25]
  wire [1:0] _T_96; // @[Cat.scala 29:58]
  wire  _T_97; // @[Shift.scala 12:21]
  wire  _T_98; // @[Shift.scala 12:21]
  wire  _T_99; // @[LZD.scala 49:16]
  wire  _T_100; // @[LZD.scala 49:27]
  wire  _T_101; // @[LZD.scala 49:25]
  wire  _T_102; // @[LZD.scala 49:47]
  wire  _T_103; // @[LZD.scala 49:59]
  wire  _T_104; // @[LZD.scala 49:35]
  wire [2:0] _T_106; // @[Cat.scala 29:58]
  wire [3:0] _T_107; // @[LZD.scala 44:32]
  wire [1:0] _T_108; // @[LZD.scala 43:32]
  wire  _T_109; // @[LZD.scala 39:14]
  wire  _T_110; // @[LZD.scala 39:21]
  wire  _T_111; // @[LZD.scala 39:30]
  wire  _T_112; // @[LZD.scala 39:27]
  wire  _T_113; // @[LZD.scala 39:25]
  wire [1:0] _T_114; // @[Cat.scala 29:58]
  wire [1:0] _T_115; // @[LZD.scala 44:32]
  wire  _T_116; // @[LZD.scala 39:14]
  wire  _T_117; // @[LZD.scala 39:21]
  wire  _T_118; // @[LZD.scala 39:30]
  wire  _T_119; // @[LZD.scala 39:27]
  wire  _T_120; // @[LZD.scala 39:25]
  wire [1:0] _T_121; // @[Cat.scala 29:58]
  wire  _T_122; // @[Shift.scala 12:21]
  wire  _T_123; // @[Shift.scala 12:21]
  wire  _T_124; // @[LZD.scala 49:16]
  wire  _T_125; // @[LZD.scala 49:27]
  wire  _T_126; // @[LZD.scala 49:25]
  wire  _T_127; // @[LZD.scala 49:47]
  wire  _T_128; // @[LZD.scala 49:59]
  wire  _T_129; // @[LZD.scala 49:35]
  wire [2:0] _T_131; // @[Cat.scala 29:58]
  wire  _T_132; // @[Shift.scala 12:21]
  wire  _T_133; // @[Shift.scala 12:21]
  wire  _T_134; // @[LZD.scala 49:16]
  wire  _T_135; // @[LZD.scala 49:27]
  wire  _T_136; // @[LZD.scala 49:25]
  wire [1:0] _T_137; // @[LZD.scala 49:47]
  wire [1:0] _T_138; // @[LZD.scala 49:59]
  wire [1:0] _T_139; // @[LZD.scala 49:35]
  wire [3:0] _T_141; // @[Cat.scala 29:58]
  wire  _T_142; // @[Shift.scala 12:21]
  wire  _T_143; // @[Shift.scala 12:21]
  wire  _T_144; // @[LZD.scala 49:16]
  wire  _T_145; // @[LZD.scala 49:27]
  wire  _T_146; // @[LZD.scala 49:25]
  wire [2:0] _T_147; // @[LZD.scala 49:47]
  wire [2:0] _T_148; // @[LZD.scala 49:59]
  wire [2:0] _T_149; // @[LZD.scala 49:35]
  wire [4:0] _T_151; // @[Cat.scala 29:58]
  wire [13:0] _T_152; // @[LZD.scala 44:32]
  wire [7:0] _T_153; // @[LZD.scala 43:32]
  wire [3:0] _T_154; // @[LZD.scala 43:32]
  wire [1:0] _T_155; // @[LZD.scala 43:32]
  wire  _T_156; // @[LZD.scala 39:14]
  wire  _T_157; // @[LZD.scala 39:21]
  wire  _T_158; // @[LZD.scala 39:30]
  wire  _T_159; // @[LZD.scala 39:27]
  wire  _T_160; // @[LZD.scala 39:25]
  wire [1:0] _T_161; // @[Cat.scala 29:58]
  wire [1:0] _T_162; // @[LZD.scala 44:32]
  wire  _T_163; // @[LZD.scala 39:14]
  wire  _T_164; // @[LZD.scala 39:21]
  wire  _T_165; // @[LZD.scala 39:30]
  wire  _T_166; // @[LZD.scala 39:27]
  wire  _T_167; // @[LZD.scala 39:25]
  wire [1:0] _T_168; // @[Cat.scala 29:58]
  wire  _T_169; // @[Shift.scala 12:21]
  wire  _T_170; // @[Shift.scala 12:21]
  wire  _T_171; // @[LZD.scala 49:16]
  wire  _T_172; // @[LZD.scala 49:27]
  wire  _T_173; // @[LZD.scala 49:25]
  wire  _T_174; // @[LZD.scala 49:47]
  wire  _T_175; // @[LZD.scala 49:59]
  wire  _T_176; // @[LZD.scala 49:35]
  wire [2:0] _T_178; // @[Cat.scala 29:58]
  wire [3:0] _T_179; // @[LZD.scala 44:32]
  wire [1:0] _T_180; // @[LZD.scala 43:32]
  wire  _T_181; // @[LZD.scala 39:14]
  wire  _T_182; // @[LZD.scala 39:21]
  wire  _T_183; // @[LZD.scala 39:30]
  wire  _T_184; // @[LZD.scala 39:27]
  wire  _T_185; // @[LZD.scala 39:25]
  wire [1:0] _T_186; // @[Cat.scala 29:58]
  wire [1:0] _T_187; // @[LZD.scala 44:32]
  wire  _T_188; // @[LZD.scala 39:14]
  wire  _T_189; // @[LZD.scala 39:21]
  wire  _T_190; // @[LZD.scala 39:30]
  wire  _T_191; // @[LZD.scala 39:27]
  wire  _T_192; // @[LZD.scala 39:25]
  wire [1:0] _T_193; // @[Cat.scala 29:58]
  wire  _T_194; // @[Shift.scala 12:21]
  wire  _T_195; // @[Shift.scala 12:21]
  wire  _T_196; // @[LZD.scala 49:16]
  wire  _T_197; // @[LZD.scala 49:27]
  wire  _T_198; // @[LZD.scala 49:25]
  wire  _T_199; // @[LZD.scala 49:47]
  wire  _T_200; // @[LZD.scala 49:59]
  wire  _T_201; // @[LZD.scala 49:35]
  wire [2:0] _T_203; // @[Cat.scala 29:58]
  wire  _T_204; // @[Shift.scala 12:21]
  wire  _T_205; // @[Shift.scala 12:21]
  wire  _T_206; // @[LZD.scala 49:16]
  wire  _T_207; // @[LZD.scala 49:27]
  wire  _T_208; // @[LZD.scala 49:25]
  wire [1:0] _T_209; // @[LZD.scala 49:47]
  wire [1:0] _T_210; // @[LZD.scala 49:59]
  wire [1:0] _T_211; // @[LZD.scala 49:35]
  wire [3:0] _T_213; // @[Cat.scala 29:58]
  wire [5:0] _T_214; // @[LZD.scala 44:32]
  wire [3:0] _T_215; // @[LZD.scala 43:32]
  wire [1:0] _T_216; // @[LZD.scala 43:32]
  wire  _T_217; // @[LZD.scala 39:14]
  wire  _T_218; // @[LZD.scala 39:21]
  wire  _T_219; // @[LZD.scala 39:30]
  wire  _T_220; // @[LZD.scala 39:27]
  wire  _T_221; // @[LZD.scala 39:25]
  wire [1:0] _T_222; // @[Cat.scala 29:58]
  wire [1:0] _T_223; // @[LZD.scala 44:32]
  wire  _T_224; // @[LZD.scala 39:14]
  wire  _T_225; // @[LZD.scala 39:21]
  wire  _T_226; // @[LZD.scala 39:30]
  wire  _T_227; // @[LZD.scala 39:27]
  wire  _T_228; // @[LZD.scala 39:25]
  wire [1:0] _T_229; // @[Cat.scala 29:58]
  wire  _T_230; // @[Shift.scala 12:21]
  wire  _T_231; // @[Shift.scala 12:21]
  wire  _T_232; // @[LZD.scala 49:16]
  wire  _T_233; // @[LZD.scala 49:27]
  wire  _T_234; // @[LZD.scala 49:25]
  wire  _T_235; // @[LZD.scala 49:47]
  wire  _T_236; // @[LZD.scala 49:59]
  wire  _T_237; // @[LZD.scala 49:35]
  wire [2:0] _T_239; // @[Cat.scala 29:58]
  wire [1:0] _T_240; // @[LZD.scala 44:32]
  wire  _T_241; // @[LZD.scala 39:14]
  wire  _T_242; // @[LZD.scala 39:21]
  wire  _T_243; // @[LZD.scala 39:30]
  wire  _T_244; // @[LZD.scala 39:27]
  wire  _T_245; // @[LZD.scala 39:25]
  wire [1:0] _T_246; // @[Cat.scala 29:58]
  wire  _T_247; // @[Shift.scala 12:21]
  wire [1:0] _T_249; // @[LZD.scala 55:32]
  wire [1:0] _T_250; // @[LZD.scala 55:20]
  wire [2:0] _T_251; // @[Cat.scala 29:58]
  wire  _T_252; // @[Shift.scala 12:21]
  wire [2:0] _T_254; // @[LZD.scala 55:32]
  wire [2:0] _T_255; // @[LZD.scala 55:20]
  wire [3:0] _T_256; // @[Cat.scala 29:58]
  wire  _T_257; // @[Shift.scala 12:21]
  wire [3:0] _T_259; // @[LZD.scala 55:32]
  wire [3:0] _T_260; // @[LZD.scala 55:20]
  wire [4:0] _T_261; // @[Cat.scala 29:58]
  wire [4:0] _T_262; // @[convert.scala 21:22]
  wire [28:0] _T_263; // @[convert.scala 22:36]
  wire  _T_264; // @[Shift.scala 16:24]
  wire  _T_266; // @[Shift.scala 12:21]
  wire [12:0] _T_267; // @[Shift.scala 64:52]
  wire [28:0] _T_269; // @[Cat.scala 29:58]
  wire [28:0] _T_270; // @[Shift.scala 64:27]
  wire [3:0] _T_271; // @[Shift.scala 66:70]
  wire  _T_272; // @[Shift.scala 12:21]
  wire [20:0] _T_273; // @[Shift.scala 64:52]
  wire [28:0] _T_275; // @[Cat.scala 29:58]
  wire [28:0] _T_276; // @[Shift.scala 64:27]
  wire [2:0] _T_277; // @[Shift.scala 66:70]
  wire  _T_278; // @[Shift.scala 12:21]
  wire [24:0] _T_279; // @[Shift.scala 64:52]
  wire [28:0] _T_281; // @[Cat.scala 29:58]
  wire [28:0] _T_282; // @[Shift.scala 64:27]
  wire [1:0] _T_283; // @[Shift.scala 66:70]
  wire  _T_284; // @[Shift.scala 12:21]
  wire [26:0] _T_285; // @[Shift.scala 64:52]
  wire [28:0] _T_287; // @[Cat.scala 29:58]
  wire [28:0] _T_288; // @[Shift.scala 64:27]
  wire  _T_289; // @[Shift.scala 66:70]
  wire [27:0] _T_291; // @[Shift.scala 64:52]
  wire [28:0] _T_292; // @[Cat.scala 29:58]
  wire [28:0] _T_293; // @[Shift.scala 64:27]
  wire [28:0] _T_294; // @[Shift.scala 16:10]
  wire  _T_295; // @[convert.scala 23:34]
  wire [27:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_297; // @[convert.scala 25:26]
  wire [4:0] _T_299; // @[convert.scala 25:42]
  wire  _T_302; // @[convert.scala 26:67]
  wire  _T_303; // @[convert.scala 26:51]
  wire [6:0] _T_304; // @[Cat.scala 29:58]
  wire [30:0] _T_306; // @[convert.scala 29:56]
  wire  _T_307; // @[convert.scala 29:60]
  wire  _T_308; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_311; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [6:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_320; // @[convert.scala 18:24]
  wire  _T_321; // @[convert.scala 18:40]
  wire  _T_322; // @[convert.scala 18:36]
  wire [29:0] _T_323; // @[convert.scala 19:24]
  wire [29:0] _T_324; // @[convert.scala 19:43]
  wire [29:0] _T_325; // @[convert.scala 19:39]
  wire [15:0] _T_326; // @[LZD.scala 43:32]
  wire [7:0] _T_327; // @[LZD.scala 43:32]
  wire [3:0] _T_328; // @[LZD.scala 43:32]
  wire [1:0] _T_329; // @[LZD.scala 43:32]
  wire  _T_330; // @[LZD.scala 39:14]
  wire  _T_331; // @[LZD.scala 39:21]
  wire  _T_332; // @[LZD.scala 39:30]
  wire  _T_333; // @[LZD.scala 39:27]
  wire  _T_334; // @[LZD.scala 39:25]
  wire [1:0] _T_335; // @[Cat.scala 29:58]
  wire [1:0] _T_336; // @[LZD.scala 44:32]
  wire  _T_337; // @[LZD.scala 39:14]
  wire  _T_338; // @[LZD.scala 39:21]
  wire  _T_339; // @[LZD.scala 39:30]
  wire  _T_340; // @[LZD.scala 39:27]
  wire  _T_341; // @[LZD.scala 39:25]
  wire [1:0] _T_342; // @[Cat.scala 29:58]
  wire  _T_343; // @[Shift.scala 12:21]
  wire  _T_344; // @[Shift.scala 12:21]
  wire  _T_345; // @[LZD.scala 49:16]
  wire  _T_346; // @[LZD.scala 49:27]
  wire  _T_347; // @[LZD.scala 49:25]
  wire  _T_348; // @[LZD.scala 49:47]
  wire  _T_349; // @[LZD.scala 49:59]
  wire  _T_350; // @[LZD.scala 49:35]
  wire [2:0] _T_352; // @[Cat.scala 29:58]
  wire [3:0] _T_353; // @[LZD.scala 44:32]
  wire [1:0] _T_354; // @[LZD.scala 43:32]
  wire  _T_355; // @[LZD.scala 39:14]
  wire  _T_356; // @[LZD.scala 39:21]
  wire  _T_357; // @[LZD.scala 39:30]
  wire  _T_358; // @[LZD.scala 39:27]
  wire  _T_359; // @[LZD.scala 39:25]
  wire [1:0] _T_360; // @[Cat.scala 29:58]
  wire [1:0] _T_361; // @[LZD.scala 44:32]
  wire  _T_362; // @[LZD.scala 39:14]
  wire  _T_363; // @[LZD.scala 39:21]
  wire  _T_364; // @[LZD.scala 39:30]
  wire  _T_365; // @[LZD.scala 39:27]
  wire  _T_366; // @[LZD.scala 39:25]
  wire [1:0] _T_367; // @[Cat.scala 29:58]
  wire  _T_368; // @[Shift.scala 12:21]
  wire  _T_369; // @[Shift.scala 12:21]
  wire  _T_370; // @[LZD.scala 49:16]
  wire  _T_371; // @[LZD.scala 49:27]
  wire  _T_372; // @[LZD.scala 49:25]
  wire  _T_373; // @[LZD.scala 49:47]
  wire  _T_374; // @[LZD.scala 49:59]
  wire  _T_375; // @[LZD.scala 49:35]
  wire [2:0] _T_377; // @[Cat.scala 29:58]
  wire  _T_378; // @[Shift.scala 12:21]
  wire  _T_379; // @[Shift.scala 12:21]
  wire  _T_380; // @[LZD.scala 49:16]
  wire  _T_381; // @[LZD.scala 49:27]
  wire  _T_382; // @[LZD.scala 49:25]
  wire [1:0] _T_383; // @[LZD.scala 49:47]
  wire [1:0] _T_384; // @[LZD.scala 49:59]
  wire [1:0] _T_385; // @[LZD.scala 49:35]
  wire [3:0] _T_387; // @[Cat.scala 29:58]
  wire [7:0] _T_388; // @[LZD.scala 44:32]
  wire [3:0] _T_389; // @[LZD.scala 43:32]
  wire [1:0] _T_390; // @[LZD.scala 43:32]
  wire  _T_391; // @[LZD.scala 39:14]
  wire  _T_392; // @[LZD.scala 39:21]
  wire  _T_393; // @[LZD.scala 39:30]
  wire  _T_394; // @[LZD.scala 39:27]
  wire  _T_395; // @[LZD.scala 39:25]
  wire [1:0] _T_396; // @[Cat.scala 29:58]
  wire [1:0] _T_397; // @[LZD.scala 44:32]
  wire  _T_398; // @[LZD.scala 39:14]
  wire  _T_399; // @[LZD.scala 39:21]
  wire  _T_400; // @[LZD.scala 39:30]
  wire  _T_401; // @[LZD.scala 39:27]
  wire  _T_402; // @[LZD.scala 39:25]
  wire [1:0] _T_403; // @[Cat.scala 29:58]
  wire  _T_404; // @[Shift.scala 12:21]
  wire  _T_405; // @[Shift.scala 12:21]
  wire  _T_406; // @[LZD.scala 49:16]
  wire  _T_407; // @[LZD.scala 49:27]
  wire  _T_408; // @[LZD.scala 49:25]
  wire  _T_409; // @[LZD.scala 49:47]
  wire  _T_410; // @[LZD.scala 49:59]
  wire  _T_411; // @[LZD.scala 49:35]
  wire [2:0] _T_413; // @[Cat.scala 29:58]
  wire [3:0] _T_414; // @[LZD.scala 44:32]
  wire [1:0] _T_415; // @[LZD.scala 43:32]
  wire  _T_416; // @[LZD.scala 39:14]
  wire  _T_417; // @[LZD.scala 39:21]
  wire  _T_418; // @[LZD.scala 39:30]
  wire  _T_419; // @[LZD.scala 39:27]
  wire  _T_420; // @[LZD.scala 39:25]
  wire [1:0] _T_421; // @[Cat.scala 29:58]
  wire [1:0] _T_422; // @[LZD.scala 44:32]
  wire  _T_423; // @[LZD.scala 39:14]
  wire  _T_424; // @[LZD.scala 39:21]
  wire  _T_425; // @[LZD.scala 39:30]
  wire  _T_426; // @[LZD.scala 39:27]
  wire  _T_427; // @[LZD.scala 39:25]
  wire [1:0] _T_428; // @[Cat.scala 29:58]
  wire  _T_429; // @[Shift.scala 12:21]
  wire  _T_430; // @[Shift.scala 12:21]
  wire  _T_431; // @[LZD.scala 49:16]
  wire  _T_432; // @[LZD.scala 49:27]
  wire  _T_433; // @[LZD.scala 49:25]
  wire  _T_434; // @[LZD.scala 49:47]
  wire  _T_435; // @[LZD.scala 49:59]
  wire  _T_436; // @[LZD.scala 49:35]
  wire [2:0] _T_438; // @[Cat.scala 29:58]
  wire  _T_439; // @[Shift.scala 12:21]
  wire  _T_440; // @[Shift.scala 12:21]
  wire  _T_441; // @[LZD.scala 49:16]
  wire  _T_442; // @[LZD.scala 49:27]
  wire  _T_443; // @[LZD.scala 49:25]
  wire [1:0] _T_444; // @[LZD.scala 49:47]
  wire [1:0] _T_445; // @[LZD.scala 49:59]
  wire [1:0] _T_446; // @[LZD.scala 49:35]
  wire [3:0] _T_448; // @[Cat.scala 29:58]
  wire  _T_449; // @[Shift.scala 12:21]
  wire  _T_450; // @[Shift.scala 12:21]
  wire  _T_451; // @[LZD.scala 49:16]
  wire  _T_452; // @[LZD.scala 49:27]
  wire  _T_453; // @[LZD.scala 49:25]
  wire [2:0] _T_454; // @[LZD.scala 49:47]
  wire [2:0] _T_455; // @[LZD.scala 49:59]
  wire [2:0] _T_456; // @[LZD.scala 49:35]
  wire [4:0] _T_458; // @[Cat.scala 29:58]
  wire [13:0] _T_459; // @[LZD.scala 44:32]
  wire [7:0] _T_460; // @[LZD.scala 43:32]
  wire [3:0] _T_461; // @[LZD.scala 43:32]
  wire [1:0] _T_462; // @[LZD.scala 43:32]
  wire  _T_463; // @[LZD.scala 39:14]
  wire  _T_464; // @[LZD.scala 39:21]
  wire  _T_465; // @[LZD.scala 39:30]
  wire  _T_466; // @[LZD.scala 39:27]
  wire  _T_467; // @[LZD.scala 39:25]
  wire [1:0] _T_468; // @[Cat.scala 29:58]
  wire [1:0] _T_469; // @[LZD.scala 44:32]
  wire  _T_470; // @[LZD.scala 39:14]
  wire  _T_471; // @[LZD.scala 39:21]
  wire  _T_472; // @[LZD.scala 39:30]
  wire  _T_473; // @[LZD.scala 39:27]
  wire  _T_474; // @[LZD.scala 39:25]
  wire [1:0] _T_475; // @[Cat.scala 29:58]
  wire  _T_476; // @[Shift.scala 12:21]
  wire  _T_477; // @[Shift.scala 12:21]
  wire  _T_478; // @[LZD.scala 49:16]
  wire  _T_479; // @[LZD.scala 49:27]
  wire  _T_480; // @[LZD.scala 49:25]
  wire  _T_481; // @[LZD.scala 49:47]
  wire  _T_482; // @[LZD.scala 49:59]
  wire  _T_483; // @[LZD.scala 49:35]
  wire [2:0] _T_485; // @[Cat.scala 29:58]
  wire [3:0] _T_486; // @[LZD.scala 44:32]
  wire [1:0] _T_487; // @[LZD.scala 43:32]
  wire  _T_488; // @[LZD.scala 39:14]
  wire  _T_489; // @[LZD.scala 39:21]
  wire  _T_490; // @[LZD.scala 39:30]
  wire  _T_491; // @[LZD.scala 39:27]
  wire  _T_492; // @[LZD.scala 39:25]
  wire [1:0] _T_493; // @[Cat.scala 29:58]
  wire [1:0] _T_494; // @[LZD.scala 44:32]
  wire  _T_495; // @[LZD.scala 39:14]
  wire  _T_496; // @[LZD.scala 39:21]
  wire  _T_497; // @[LZD.scala 39:30]
  wire  _T_498; // @[LZD.scala 39:27]
  wire  _T_499; // @[LZD.scala 39:25]
  wire [1:0] _T_500; // @[Cat.scala 29:58]
  wire  _T_501; // @[Shift.scala 12:21]
  wire  _T_502; // @[Shift.scala 12:21]
  wire  _T_503; // @[LZD.scala 49:16]
  wire  _T_504; // @[LZD.scala 49:27]
  wire  _T_505; // @[LZD.scala 49:25]
  wire  _T_506; // @[LZD.scala 49:47]
  wire  _T_507; // @[LZD.scala 49:59]
  wire  _T_508; // @[LZD.scala 49:35]
  wire [2:0] _T_510; // @[Cat.scala 29:58]
  wire  _T_511; // @[Shift.scala 12:21]
  wire  _T_512; // @[Shift.scala 12:21]
  wire  _T_513; // @[LZD.scala 49:16]
  wire  _T_514; // @[LZD.scala 49:27]
  wire  _T_515; // @[LZD.scala 49:25]
  wire [1:0] _T_516; // @[LZD.scala 49:47]
  wire [1:0] _T_517; // @[LZD.scala 49:59]
  wire [1:0] _T_518; // @[LZD.scala 49:35]
  wire [3:0] _T_520; // @[Cat.scala 29:58]
  wire [5:0] _T_521; // @[LZD.scala 44:32]
  wire [3:0] _T_522; // @[LZD.scala 43:32]
  wire [1:0] _T_523; // @[LZD.scala 43:32]
  wire  _T_524; // @[LZD.scala 39:14]
  wire  _T_525; // @[LZD.scala 39:21]
  wire  _T_526; // @[LZD.scala 39:30]
  wire  _T_527; // @[LZD.scala 39:27]
  wire  _T_528; // @[LZD.scala 39:25]
  wire [1:0] _T_529; // @[Cat.scala 29:58]
  wire [1:0] _T_530; // @[LZD.scala 44:32]
  wire  _T_531; // @[LZD.scala 39:14]
  wire  _T_532; // @[LZD.scala 39:21]
  wire  _T_533; // @[LZD.scala 39:30]
  wire  _T_534; // @[LZD.scala 39:27]
  wire  _T_535; // @[LZD.scala 39:25]
  wire [1:0] _T_536; // @[Cat.scala 29:58]
  wire  _T_537; // @[Shift.scala 12:21]
  wire  _T_538; // @[Shift.scala 12:21]
  wire  _T_539; // @[LZD.scala 49:16]
  wire  _T_540; // @[LZD.scala 49:27]
  wire  _T_541; // @[LZD.scala 49:25]
  wire  _T_542; // @[LZD.scala 49:47]
  wire  _T_543; // @[LZD.scala 49:59]
  wire  _T_544; // @[LZD.scala 49:35]
  wire [2:0] _T_546; // @[Cat.scala 29:58]
  wire [1:0] _T_547; // @[LZD.scala 44:32]
  wire  _T_548; // @[LZD.scala 39:14]
  wire  _T_549; // @[LZD.scala 39:21]
  wire  _T_550; // @[LZD.scala 39:30]
  wire  _T_551; // @[LZD.scala 39:27]
  wire  _T_552; // @[LZD.scala 39:25]
  wire [1:0] _T_553; // @[Cat.scala 29:58]
  wire  _T_554; // @[Shift.scala 12:21]
  wire [1:0] _T_556; // @[LZD.scala 55:32]
  wire [1:0] _T_557; // @[LZD.scala 55:20]
  wire [2:0] _T_558; // @[Cat.scala 29:58]
  wire  _T_559; // @[Shift.scala 12:21]
  wire [2:0] _T_561; // @[LZD.scala 55:32]
  wire [2:0] _T_562; // @[LZD.scala 55:20]
  wire [3:0] _T_563; // @[Cat.scala 29:58]
  wire  _T_564; // @[Shift.scala 12:21]
  wire [3:0] _T_566; // @[LZD.scala 55:32]
  wire [3:0] _T_567; // @[LZD.scala 55:20]
  wire [4:0] _T_568; // @[Cat.scala 29:58]
  wire [4:0] _T_569; // @[convert.scala 21:22]
  wire [28:0] _T_570; // @[convert.scala 22:36]
  wire  _T_571; // @[Shift.scala 16:24]
  wire  _T_573; // @[Shift.scala 12:21]
  wire [12:0] _T_574; // @[Shift.scala 64:52]
  wire [28:0] _T_576; // @[Cat.scala 29:58]
  wire [28:0] _T_577; // @[Shift.scala 64:27]
  wire [3:0] _T_578; // @[Shift.scala 66:70]
  wire  _T_579; // @[Shift.scala 12:21]
  wire [20:0] _T_580; // @[Shift.scala 64:52]
  wire [28:0] _T_582; // @[Cat.scala 29:58]
  wire [28:0] _T_583; // @[Shift.scala 64:27]
  wire [2:0] _T_584; // @[Shift.scala 66:70]
  wire  _T_585; // @[Shift.scala 12:21]
  wire [24:0] _T_586; // @[Shift.scala 64:52]
  wire [28:0] _T_588; // @[Cat.scala 29:58]
  wire [28:0] _T_589; // @[Shift.scala 64:27]
  wire [1:0] _T_590; // @[Shift.scala 66:70]
  wire  _T_591; // @[Shift.scala 12:21]
  wire [26:0] _T_592; // @[Shift.scala 64:52]
  wire [28:0] _T_594; // @[Cat.scala 29:58]
  wire [28:0] _T_595; // @[Shift.scala 64:27]
  wire  _T_596; // @[Shift.scala 66:70]
  wire [27:0] _T_598; // @[Shift.scala 64:52]
  wire [28:0] _T_599; // @[Cat.scala 29:58]
  wire [28:0] _T_600; // @[Shift.scala 64:27]
  wire [28:0] _T_601; // @[Shift.scala 16:10]
  wire  _T_602; // @[convert.scala 23:34]
  wire [27:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_604; // @[convert.scala 25:26]
  wire [4:0] _T_606; // @[convert.scala 25:42]
  wire  _T_609; // @[convert.scala 26:67]
  wire  _T_610; // @[convert.scala 26:51]
  wire [6:0] _T_611; // @[Cat.scala 29:58]
  wire [30:0] _T_613; // @[convert.scala 29:56]
  wire  _T_614; // @[convert.scala 29:60]
  wire  _T_615; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_618; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [6:0] decB_scale; // @[convert.scala 32:24]
  wire  _T_627; // @[convert.scala 18:24]
  wire  _T_628; // @[convert.scala 18:40]
  wire  _T_629; // @[convert.scala 18:36]
  wire [29:0] _T_630; // @[convert.scala 19:24]
  wire [29:0] _T_631; // @[convert.scala 19:43]
  wire [29:0] _T_632; // @[convert.scala 19:39]
  wire [15:0] _T_633; // @[LZD.scala 43:32]
  wire [7:0] _T_634; // @[LZD.scala 43:32]
  wire [3:0] _T_635; // @[LZD.scala 43:32]
  wire [1:0] _T_636; // @[LZD.scala 43:32]
  wire  _T_637; // @[LZD.scala 39:14]
  wire  _T_638; // @[LZD.scala 39:21]
  wire  _T_639; // @[LZD.scala 39:30]
  wire  _T_640; // @[LZD.scala 39:27]
  wire  _T_641; // @[LZD.scala 39:25]
  wire [1:0] _T_642; // @[Cat.scala 29:58]
  wire [1:0] _T_643; // @[LZD.scala 44:32]
  wire  _T_644; // @[LZD.scala 39:14]
  wire  _T_645; // @[LZD.scala 39:21]
  wire  _T_646; // @[LZD.scala 39:30]
  wire  _T_647; // @[LZD.scala 39:27]
  wire  _T_648; // @[LZD.scala 39:25]
  wire [1:0] _T_649; // @[Cat.scala 29:58]
  wire  _T_650; // @[Shift.scala 12:21]
  wire  _T_651; // @[Shift.scala 12:21]
  wire  _T_652; // @[LZD.scala 49:16]
  wire  _T_653; // @[LZD.scala 49:27]
  wire  _T_654; // @[LZD.scala 49:25]
  wire  _T_655; // @[LZD.scala 49:47]
  wire  _T_656; // @[LZD.scala 49:59]
  wire  _T_657; // @[LZD.scala 49:35]
  wire [2:0] _T_659; // @[Cat.scala 29:58]
  wire [3:0] _T_660; // @[LZD.scala 44:32]
  wire [1:0] _T_661; // @[LZD.scala 43:32]
  wire  _T_662; // @[LZD.scala 39:14]
  wire  _T_663; // @[LZD.scala 39:21]
  wire  _T_664; // @[LZD.scala 39:30]
  wire  _T_665; // @[LZD.scala 39:27]
  wire  _T_666; // @[LZD.scala 39:25]
  wire [1:0] _T_667; // @[Cat.scala 29:58]
  wire [1:0] _T_668; // @[LZD.scala 44:32]
  wire  _T_669; // @[LZD.scala 39:14]
  wire  _T_670; // @[LZD.scala 39:21]
  wire  _T_671; // @[LZD.scala 39:30]
  wire  _T_672; // @[LZD.scala 39:27]
  wire  _T_673; // @[LZD.scala 39:25]
  wire [1:0] _T_674; // @[Cat.scala 29:58]
  wire  _T_675; // @[Shift.scala 12:21]
  wire  _T_676; // @[Shift.scala 12:21]
  wire  _T_677; // @[LZD.scala 49:16]
  wire  _T_678; // @[LZD.scala 49:27]
  wire  _T_679; // @[LZD.scala 49:25]
  wire  _T_680; // @[LZD.scala 49:47]
  wire  _T_681; // @[LZD.scala 49:59]
  wire  _T_682; // @[LZD.scala 49:35]
  wire [2:0] _T_684; // @[Cat.scala 29:58]
  wire  _T_685; // @[Shift.scala 12:21]
  wire  _T_686; // @[Shift.scala 12:21]
  wire  _T_687; // @[LZD.scala 49:16]
  wire  _T_688; // @[LZD.scala 49:27]
  wire  _T_689; // @[LZD.scala 49:25]
  wire [1:0] _T_690; // @[LZD.scala 49:47]
  wire [1:0] _T_691; // @[LZD.scala 49:59]
  wire [1:0] _T_692; // @[LZD.scala 49:35]
  wire [3:0] _T_694; // @[Cat.scala 29:58]
  wire [7:0] _T_695; // @[LZD.scala 44:32]
  wire [3:0] _T_696; // @[LZD.scala 43:32]
  wire [1:0] _T_697; // @[LZD.scala 43:32]
  wire  _T_698; // @[LZD.scala 39:14]
  wire  _T_699; // @[LZD.scala 39:21]
  wire  _T_700; // @[LZD.scala 39:30]
  wire  _T_701; // @[LZD.scala 39:27]
  wire  _T_702; // @[LZD.scala 39:25]
  wire [1:0] _T_703; // @[Cat.scala 29:58]
  wire [1:0] _T_704; // @[LZD.scala 44:32]
  wire  _T_705; // @[LZD.scala 39:14]
  wire  _T_706; // @[LZD.scala 39:21]
  wire  _T_707; // @[LZD.scala 39:30]
  wire  _T_708; // @[LZD.scala 39:27]
  wire  _T_709; // @[LZD.scala 39:25]
  wire [1:0] _T_710; // @[Cat.scala 29:58]
  wire  _T_711; // @[Shift.scala 12:21]
  wire  _T_712; // @[Shift.scala 12:21]
  wire  _T_713; // @[LZD.scala 49:16]
  wire  _T_714; // @[LZD.scala 49:27]
  wire  _T_715; // @[LZD.scala 49:25]
  wire  _T_716; // @[LZD.scala 49:47]
  wire  _T_717; // @[LZD.scala 49:59]
  wire  _T_718; // @[LZD.scala 49:35]
  wire [2:0] _T_720; // @[Cat.scala 29:58]
  wire [3:0] _T_721; // @[LZD.scala 44:32]
  wire [1:0] _T_722; // @[LZD.scala 43:32]
  wire  _T_723; // @[LZD.scala 39:14]
  wire  _T_724; // @[LZD.scala 39:21]
  wire  _T_725; // @[LZD.scala 39:30]
  wire  _T_726; // @[LZD.scala 39:27]
  wire  _T_727; // @[LZD.scala 39:25]
  wire [1:0] _T_728; // @[Cat.scala 29:58]
  wire [1:0] _T_729; // @[LZD.scala 44:32]
  wire  _T_730; // @[LZD.scala 39:14]
  wire  _T_731; // @[LZD.scala 39:21]
  wire  _T_732; // @[LZD.scala 39:30]
  wire  _T_733; // @[LZD.scala 39:27]
  wire  _T_734; // @[LZD.scala 39:25]
  wire [1:0] _T_735; // @[Cat.scala 29:58]
  wire  _T_736; // @[Shift.scala 12:21]
  wire  _T_737; // @[Shift.scala 12:21]
  wire  _T_738; // @[LZD.scala 49:16]
  wire  _T_739; // @[LZD.scala 49:27]
  wire  _T_740; // @[LZD.scala 49:25]
  wire  _T_741; // @[LZD.scala 49:47]
  wire  _T_742; // @[LZD.scala 49:59]
  wire  _T_743; // @[LZD.scala 49:35]
  wire [2:0] _T_745; // @[Cat.scala 29:58]
  wire  _T_746; // @[Shift.scala 12:21]
  wire  _T_747; // @[Shift.scala 12:21]
  wire  _T_748; // @[LZD.scala 49:16]
  wire  _T_749; // @[LZD.scala 49:27]
  wire  _T_750; // @[LZD.scala 49:25]
  wire [1:0] _T_751; // @[LZD.scala 49:47]
  wire [1:0] _T_752; // @[LZD.scala 49:59]
  wire [1:0] _T_753; // @[LZD.scala 49:35]
  wire [3:0] _T_755; // @[Cat.scala 29:58]
  wire  _T_756; // @[Shift.scala 12:21]
  wire  _T_757; // @[Shift.scala 12:21]
  wire  _T_758; // @[LZD.scala 49:16]
  wire  _T_759; // @[LZD.scala 49:27]
  wire  _T_760; // @[LZD.scala 49:25]
  wire [2:0] _T_761; // @[LZD.scala 49:47]
  wire [2:0] _T_762; // @[LZD.scala 49:59]
  wire [2:0] _T_763; // @[LZD.scala 49:35]
  wire [4:0] _T_765; // @[Cat.scala 29:58]
  wire [13:0] _T_766; // @[LZD.scala 44:32]
  wire [7:0] _T_767; // @[LZD.scala 43:32]
  wire [3:0] _T_768; // @[LZD.scala 43:32]
  wire [1:0] _T_769; // @[LZD.scala 43:32]
  wire  _T_770; // @[LZD.scala 39:14]
  wire  _T_771; // @[LZD.scala 39:21]
  wire  _T_772; // @[LZD.scala 39:30]
  wire  _T_773; // @[LZD.scala 39:27]
  wire  _T_774; // @[LZD.scala 39:25]
  wire [1:0] _T_775; // @[Cat.scala 29:58]
  wire [1:0] _T_776; // @[LZD.scala 44:32]
  wire  _T_777; // @[LZD.scala 39:14]
  wire  _T_778; // @[LZD.scala 39:21]
  wire  _T_779; // @[LZD.scala 39:30]
  wire  _T_780; // @[LZD.scala 39:27]
  wire  _T_781; // @[LZD.scala 39:25]
  wire [1:0] _T_782; // @[Cat.scala 29:58]
  wire  _T_783; // @[Shift.scala 12:21]
  wire  _T_784; // @[Shift.scala 12:21]
  wire  _T_785; // @[LZD.scala 49:16]
  wire  _T_786; // @[LZD.scala 49:27]
  wire  _T_787; // @[LZD.scala 49:25]
  wire  _T_788; // @[LZD.scala 49:47]
  wire  _T_789; // @[LZD.scala 49:59]
  wire  _T_790; // @[LZD.scala 49:35]
  wire [2:0] _T_792; // @[Cat.scala 29:58]
  wire [3:0] _T_793; // @[LZD.scala 44:32]
  wire [1:0] _T_794; // @[LZD.scala 43:32]
  wire  _T_795; // @[LZD.scala 39:14]
  wire  _T_796; // @[LZD.scala 39:21]
  wire  _T_797; // @[LZD.scala 39:30]
  wire  _T_798; // @[LZD.scala 39:27]
  wire  _T_799; // @[LZD.scala 39:25]
  wire [1:0] _T_800; // @[Cat.scala 29:58]
  wire [1:0] _T_801; // @[LZD.scala 44:32]
  wire  _T_802; // @[LZD.scala 39:14]
  wire  _T_803; // @[LZD.scala 39:21]
  wire  _T_804; // @[LZD.scala 39:30]
  wire  _T_805; // @[LZD.scala 39:27]
  wire  _T_806; // @[LZD.scala 39:25]
  wire [1:0] _T_807; // @[Cat.scala 29:58]
  wire  _T_808; // @[Shift.scala 12:21]
  wire  _T_809; // @[Shift.scala 12:21]
  wire  _T_810; // @[LZD.scala 49:16]
  wire  _T_811; // @[LZD.scala 49:27]
  wire  _T_812; // @[LZD.scala 49:25]
  wire  _T_813; // @[LZD.scala 49:47]
  wire  _T_814; // @[LZD.scala 49:59]
  wire  _T_815; // @[LZD.scala 49:35]
  wire [2:0] _T_817; // @[Cat.scala 29:58]
  wire  _T_818; // @[Shift.scala 12:21]
  wire  _T_819; // @[Shift.scala 12:21]
  wire  _T_820; // @[LZD.scala 49:16]
  wire  _T_821; // @[LZD.scala 49:27]
  wire  _T_822; // @[LZD.scala 49:25]
  wire [1:0] _T_823; // @[LZD.scala 49:47]
  wire [1:0] _T_824; // @[LZD.scala 49:59]
  wire [1:0] _T_825; // @[LZD.scala 49:35]
  wire [3:0] _T_827; // @[Cat.scala 29:58]
  wire [5:0] _T_828; // @[LZD.scala 44:32]
  wire [3:0] _T_829; // @[LZD.scala 43:32]
  wire [1:0] _T_830; // @[LZD.scala 43:32]
  wire  _T_831; // @[LZD.scala 39:14]
  wire  _T_832; // @[LZD.scala 39:21]
  wire  _T_833; // @[LZD.scala 39:30]
  wire  _T_834; // @[LZD.scala 39:27]
  wire  _T_835; // @[LZD.scala 39:25]
  wire [1:0] _T_836; // @[Cat.scala 29:58]
  wire [1:0] _T_837; // @[LZD.scala 44:32]
  wire  _T_838; // @[LZD.scala 39:14]
  wire  _T_839; // @[LZD.scala 39:21]
  wire  _T_840; // @[LZD.scala 39:30]
  wire  _T_841; // @[LZD.scala 39:27]
  wire  _T_842; // @[LZD.scala 39:25]
  wire [1:0] _T_843; // @[Cat.scala 29:58]
  wire  _T_844; // @[Shift.scala 12:21]
  wire  _T_845; // @[Shift.scala 12:21]
  wire  _T_846; // @[LZD.scala 49:16]
  wire  _T_847; // @[LZD.scala 49:27]
  wire  _T_848; // @[LZD.scala 49:25]
  wire  _T_849; // @[LZD.scala 49:47]
  wire  _T_850; // @[LZD.scala 49:59]
  wire  _T_851; // @[LZD.scala 49:35]
  wire [2:0] _T_853; // @[Cat.scala 29:58]
  wire [1:0] _T_854; // @[LZD.scala 44:32]
  wire  _T_855; // @[LZD.scala 39:14]
  wire  _T_856; // @[LZD.scala 39:21]
  wire  _T_857; // @[LZD.scala 39:30]
  wire  _T_858; // @[LZD.scala 39:27]
  wire  _T_859; // @[LZD.scala 39:25]
  wire [1:0] _T_860; // @[Cat.scala 29:58]
  wire  _T_861; // @[Shift.scala 12:21]
  wire [1:0] _T_863; // @[LZD.scala 55:32]
  wire [1:0] _T_864; // @[LZD.scala 55:20]
  wire [2:0] _T_865; // @[Cat.scala 29:58]
  wire  _T_866; // @[Shift.scala 12:21]
  wire [2:0] _T_868; // @[LZD.scala 55:32]
  wire [2:0] _T_869; // @[LZD.scala 55:20]
  wire [3:0] _T_870; // @[Cat.scala 29:58]
  wire  _T_871; // @[Shift.scala 12:21]
  wire [3:0] _T_873; // @[LZD.scala 55:32]
  wire [3:0] _T_874; // @[LZD.scala 55:20]
  wire [4:0] _T_875; // @[Cat.scala 29:58]
  wire [4:0] _T_876; // @[convert.scala 21:22]
  wire [28:0] _T_877; // @[convert.scala 22:36]
  wire  _T_878; // @[Shift.scala 16:24]
  wire  _T_880; // @[Shift.scala 12:21]
  wire [12:0] _T_881; // @[Shift.scala 64:52]
  wire [28:0] _T_883; // @[Cat.scala 29:58]
  wire [28:0] _T_884; // @[Shift.scala 64:27]
  wire [3:0] _T_885; // @[Shift.scala 66:70]
  wire  _T_886; // @[Shift.scala 12:21]
  wire [20:0] _T_887; // @[Shift.scala 64:52]
  wire [28:0] _T_889; // @[Cat.scala 29:58]
  wire [28:0] _T_890; // @[Shift.scala 64:27]
  wire [2:0] _T_891; // @[Shift.scala 66:70]
  wire  _T_892; // @[Shift.scala 12:21]
  wire [24:0] _T_893; // @[Shift.scala 64:52]
  wire [28:0] _T_895; // @[Cat.scala 29:58]
  wire [28:0] _T_896; // @[Shift.scala 64:27]
  wire [1:0] _T_897; // @[Shift.scala 66:70]
  wire  _T_898; // @[Shift.scala 12:21]
  wire [26:0] _T_899; // @[Shift.scala 64:52]
  wire [28:0] _T_901; // @[Cat.scala 29:58]
  wire [28:0] _T_902; // @[Shift.scala 64:27]
  wire  _T_903; // @[Shift.scala 66:70]
  wire [27:0] _T_905; // @[Shift.scala 64:52]
  wire [28:0] _T_906; // @[Cat.scala 29:58]
  wire [28:0] _T_907; // @[Shift.scala 64:27]
  wire [28:0] _T_908; // @[Shift.scala 16:10]
  wire  _T_909; // @[convert.scala 23:34]
  wire [27:0] decC_fraction; // @[convert.scala 24:34]
  wire  _T_911; // @[convert.scala 25:26]
  wire [4:0] _T_913; // @[convert.scala 25:42]
  wire  _T_916; // @[convert.scala 26:67]
  wire  _T_917; // @[convert.scala 26:51]
  wire [6:0] _T_918; // @[Cat.scala 29:58]
  wire [30:0] _T_920; // @[convert.scala 29:56]
  wire  _T_921; // @[convert.scala 29:60]
  wire  _T_922; // @[convert.scala 29:41]
  wire  decC_isNaR; // @[convert.scala 29:39]
  wire  _T_925; // @[convert.scala 30:19]
  wire  decC_isZero; // @[convert.scala 30:41]
  wire [6:0] decC_scale; // @[convert.scala 32:24]
  wire  _T_933; // @[PositFMA.scala 58:30]
  wire  outIsNaR; // @[PositFMA.scala 58:44]
  wire  _T_934; // @[PositFMA.scala 59:34]
  wire  _T_935; // @[PositFMA.scala 59:47]
  wire  _T_936; // @[PositFMA.scala 59:45]
  wire [29:0] _T_938; // @[Cat.scala 29:58]
  wire [29:0] sigA; // @[PositFMA.scala 59:76]
  wire  _T_939; // @[PositFMA.scala 60:34]
  wire  _T_940; // @[PositFMA.scala 60:47]
  wire  _T_941; // @[PositFMA.scala 60:45]
  wire [29:0] _T_943; // @[Cat.scala 29:58]
  wire [29:0] sigB; // @[PositFMA.scala 60:76]
  wire [59:0] _T_944; // @[PositFMA.scala 61:25]
  wire [59:0] sigP; // @[PositFMA.scala 61:33]
  wire [1:0] head2; // @[PositFMA.scala 62:28]
  wire  _T_945; // @[PositFMA.scala 63:31]
  wire  _T_946; // @[PositFMA.scala 63:25]
  wire  _T_947; // @[PositFMA.scala 63:42]
  wire  addTwo; // @[PositFMA.scala 63:35]
  wire  _T_948; // @[PositFMA.scala 65:23]
  wire  _T_949; // @[PositFMA.scala 65:49]
  wire  addOne; // @[PositFMA.scala 65:43]
  wire [1:0] _T_950; // @[Cat.scala 29:58]
  wire [2:0] expBias; // @[PositFMA.scala 66:39]
  wire  mulSign; // @[PositFMA.scala 67:28]
  wire [7:0] _T_951; // @[PositFMA.scala 69:30]
  wire [7:0] _GEN_12; // @[PositFMA.scala 69:44]
  wire [7:0] _T_953; // @[PositFMA.scala 69:44]
  wire [7:0] mulScale; // @[PositFMA.scala 69:44]
  wire [57:0] _T_954; // @[PositFMA.scala 72:29]
  wire [56:0] _T_955; // @[PositFMA.scala 73:29]
  wire [57:0] _T_956; // @[PositFMA.scala 73:48]
  wire [57:0] mulSigTmp; // @[PositFMA.scala 70:22]
  wire  _T_958; // @[PositFMA.scala 77:39]
  wire  _T_959; // @[PositFMA.scala 77:43]
  wire [56:0] _T_960; // @[PositFMA.scala 78:39]
  wire [58:0] mulSig; // @[Cat.scala 29:58]
  reg  outIsNaR_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg [58:0] mulSig_phase2; // @[Reg.scala 15:16]
  reg [63:0] _RAND_1;
  reg [27:0] addFrac_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [7:0] mulScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [6:0] addScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  addSign_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  addZero_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  inValid_phase2; // @[Valid.scala 117:22]
  reg [31:0] _RAND_7;
  wire  _T_986; // @[PositFMA.scala 107:29]
  wire  _T_987; // @[PositFMA.scala 107:47]
  wire  _T_988; // @[PositFMA.scala 107:45]
  wire [58:0] extAddSig; // @[Cat.scala 29:58]
  wire [7:0] _GEN_13; // @[PositFMA.scala 111:39]
  wire  mulGreater; // @[PositFMA.scala 111:39]
  wire [7:0] greaterScale; // @[PositFMA.scala 112:26]
  wire [7:0] smallerScale; // @[PositFMA.scala 113:26]
  wire [7:0] _T_992; // @[PositFMA.scala 114:36]
  wire [7:0] scaleDiff; // @[PositFMA.scala 114:36]
  wire [58:0] greaterSig; // @[PositFMA.scala 115:26]
  wire [58:0] smallerSigTmp; // @[PositFMA.scala 116:26]
  wire [7:0] _T_993; // @[PositFMA.scala 117:69]
  wire  _T_994; // @[Shift.scala 39:24]
  wire [5:0] _T_995; // @[Shift.scala 40:44]
  wire [26:0] _T_996; // @[Shift.scala 90:30]
  wire [31:0] _T_997; // @[Shift.scala 90:48]
  wire  _T_998; // @[Shift.scala 90:57]
  wire [26:0] _GEN_14; // @[Shift.scala 90:39]
  wire [26:0] _T_999; // @[Shift.scala 90:39]
  wire  _T_1000; // @[Shift.scala 12:21]
  wire  _T_1001; // @[Shift.scala 12:21]
  wire [31:0] _T_1003; // @[Bitwise.scala 71:12]
  wire [58:0] _T_1004; // @[Cat.scala 29:58]
  wire [58:0] _T_1005; // @[Shift.scala 91:22]
  wire [4:0] _T_1006; // @[Shift.scala 92:77]
  wire [42:0] _T_1007; // @[Shift.scala 90:30]
  wire [15:0] _T_1008; // @[Shift.scala 90:48]
  wire  _T_1009; // @[Shift.scala 90:57]
  wire [42:0] _GEN_15; // @[Shift.scala 90:39]
  wire [42:0] _T_1010; // @[Shift.scala 90:39]
  wire  _T_1011; // @[Shift.scala 12:21]
  wire  _T_1012; // @[Shift.scala 12:21]
  wire [15:0] _T_1014; // @[Bitwise.scala 71:12]
  wire [58:0] _T_1015; // @[Cat.scala 29:58]
  wire [58:0] _T_1016; // @[Shift.scala 91:22]
  wire [3:0] _T_1017; // @[Shift.scala 92:77]
  wire [50:0] _T_1018; // @[Shift.scala 90:30]
  wire [7:0] _T_1019; // @[Shift.scala 90:48]
  wire  _T_1020; // @[Shift.scala 90:57]
  wire [50:0] _GEN_16; // @[Shift.scala 90:39]
  wire [50:0] _T_1021; // @[Shift.scala 90:39]
  wire  _T_1022; // @[Shift.scala 12:21]
  wire  _T_1023; // @[Shift.scala 12:21]
  wire [7:0] _T_1025; // @[Bitwise.scala 71:12]
  wire [58:0] _T_1026; // @[Cat.scala 29:58]
  wire [58:0] _T_1027; // @[Shift.scala 91:22]
  wire [2:0] _T_1028; // @[Shift.scala 92:77]
  wire [54:0] _T_1029; // @[Shift.scala 90:30]
  wire [3:0] _T_1030; // @[Shift.scala 90:48]
  wire  _T_1031; // @[Shift.scala 90:57]
  wire [54:0] _GEN_17; // @[Shift.scala 90:39]
  wire [54:0] _T_1032; // @[Shift.scala 90:39]
  wire  _T_1033; // @[Shift.scala 12:21]
  wire  _T_1034; // @[Shift.scala 12:21]
  wire [3:0] _T_1036; // @[Bitwise.scala 71:12]
  wire [58:0] _T_1037; // @[Cat.scala 29:58]
  wire [58:0] _T_1038; // @[Shift.scala 91:22]
  wire [1:0] _T_1039; // @[Shift.scala 92:77]
  wire [56:0] _T_1040; // @[Shift.scala 90:30]
  wire [1:0] _T_1041; // @[Shift.scala 90:48]
  wire  _T_1042; // @[Shift.scala 90:57]
  wire [56:0] _GEN_18; // @[Shift.scala 90:39]
  wire [56:0] _T_1043; // @[Shift.scala 90:39]
  wire  _T_1044; // @[Shift.scala 12:21]
  wire  _T_1045; // @[Shift.scala 12:21]
  wire [1:0] _T_1047; // @[Bitwise.scala 71:12]
  wire [58:0] _T_1048; // @[Cat.scala 29:58]
  wire [58:0] _T_1049; // @[Shift.scala 91:22]
  wire  _T_1050; // @[Shift.scala 92:77]
  wire [57:0] _T_1051; // @[Shift.scala 90:30]
  wire  _T_1052; // @[Shift.scala 90:48]
  wire [57:0] _GEN_19; // @[Shift.scala 90:39]
  wire [57:0] _T_1054; // @[Shift.scala 90:39]
  wire  _T_1056; // @[Shift.scala 12:21]
  wire [58:0] _T_1057; // @[Cat.scala 29:58]
  wire [58:0] _T_1058; // @[Shift.scala 91:22]
  wire [58:0] _T_1061; // @[Bitwise.scala 71:12]
  wire [58:0] smallerSig; // @[Shift.scala 39:10]
  wire [59:0] rawSumSig; // @[PositFMA.scala 118:34]
  wire  _T_1062; // @[PositFMA.scala 119:42]
  wire  _T_1063; // @[PositFMA.scala 119:46]
  wire  _T_1064; // @[PositFMA.scala 119:79]
  wire  sumSign; // @[PositFMA.scala 119:63]
  wire [58:0] _T_1066; // @[PositFMA.scala 120:50]
  wire [59:0] signSumSig; // @[Cat.scala 29:58]
  wire [58:0] _T_1067; // @[PositFMA.scala 124:33]
  wire [58:0] _T_1068; // @[PositFMA.scala 124:68]
  wire [58:0] sumXor; // @[PositFMA.scala 124:51]
  wire [31:0] _T_1069; // @[LZD.scala 43:32]
  wire [15:0] _T_1070; // @[LZD.scala 43:32]
  wire [7:0] _T_1071; // @[LZD.scala 43:32]
  wire [3:0] _T_1072; // @[LZD.scala 43:32]
  wire [1:0] _T_1073; // @[LZD.scala 43:32]
  wire  _T_1074; // @[LZD.scala 39:14]
  wire  _T_1075; // @[LZD.scala 39:21]
  wire  _T_1076; // @[LZD.scala 39:30]
  wire  _T_1077; // @[LZD.scala 39:27]
  wire  _T_1078; // @[LZD.scala 39:25]
  wire [1:0] _T_1079; // @[Cat.scala 29:58]
  wire [1:0] _T_1080; // @[LZD.scala 44:32]
  wire  _T_1081; // @[LZD.scala 39:14]
  wire  _T_1082; // @[LZD.scala 39:21]
  wire  _T_1083; // @[LZD.scala 39:30]
  wire  _T_1084; // @[LZD.scala 39:27]
  wire  _T_1085; // @[LZD.scala 39:25]
  wire [1:0] _T_1086; // @[Cat.scala 29:58]
  wire  _T_1087; // @[Shift.scala 12:21]
  wire  _T_1088; // @[Shift.scala 12:21]
  wire  _T_1089; // @[LZD.scala 49:16]
  wire  _T_1090; // @[LZD.scala 49:27]
  wire  _T_1091; // @[LZD.scala 49:25]
  wire  _T_1092; // @[LZD.scala 49:47]
  wire  _T_1093; // @[LZD.scala 49:59]
  wire  _T_1094; // @[LZD.scala 49:35]
  wire [2:0] _T_1096; // @[Cat.scala 29:58]
  wire [3:0] _T_1097; // @[LZD.scala 44:32]
  wire [1:0] _T_1098; // @[LZD.scala 43:32]
  wire  _T_1099; // @[LZD.scala 39:14]
  wire  _T_1100; // @[LZD.scala 39:21]
  wire  _T_1101; // @[LZD.scala 39:30]
  wire  _T_1102; // @[LZD.scala 39:27]
  wire  _T_1103; // @[LZD.scala 39:25]
  wire [1:0] _T_1104; // @[Cat.scala 29:58]
  wire [1:0] _T_1105; // @[LZD.scala 44:32]
  wire  _T_1106; // @[LZD.scala 39:14]
  wire  _T_1107; // @[LZD.scala 39:21]
  wire  _T_1108; // @[LZD.scala 39:30]
  wire  _T_1109; // @[LZD.scala 39:27]
  wire  _T_1110; // @[LZD.scala 39:25]
  wire [1:0] _T_1111; // @[Cat.scala 29:58]
  wire  _T_1112; // @[Shift.scala 12:21]
  wire  _T_1113; // @[Shift.scala 12:21]
  wire  _T_1114; // @[LZD.scala 49:16]
  wire  _T_1115; // @[LZD.scala 49:27]
  wire  _T_1116; // @[LZD.scala 49:25]
  wire  _T_1117; // @[LZD.scala 49:47]
  wire  _T_1118; // @[LZD.scala 49:59]
  wire  _T_1119; // @[LZD.scala 49:35]
  wire [2:0] _T_1121; // @[Cat.scala 29:58]
  wire  _T_1122; // @[Shift.scala 12:21]
  wire  _T_1123; // @[Shift.scala 12:21]
  wire  _T_1124; // @[LZD.scala 49:16]
  wire  _T_1125; // @[LZD.scala 49:27]
  wire  _T_1126; // @[LZD.scala 49:25]
  wire [1:0] _T_1127; // @[LZD.scala 49:47]
  wire [1:0] _T_1128; // @[LZD.scala 49:59]
  wire [1:0] _T_1129; // @[LZD.scala 49:35]
  wire [3:0] _T_1131; // @[Cat.scala 29:58]
  wire [7:0] _T_1132; // @[LZD.scala 44:32]
  wire [3:0] _T_1133; // @[LZD.scala 43:32]
  wire [1:0] _T_1134; // @[LZD.scala 43:32]
  wire  _T_1135; // @[LZD.scala 39:14]
  wire  _T_1136; // @[LZD.scala 39:21]
  wire  _T_1137; // @[LZD.scala 39:30]
  wire  _T_1138; // @[LZD.scala 39:27]
  wire  _T_1139; // @[LZD.scala 39:25]
  wire [1:0] _T_1140; // @[Cat.scala 29:58]
  wire [1:0] _T_1141; // @[LZD.scala 44:32]
  wire  _T_1142; // @[LZD.scala 39:14]
  wire  _T_1143; // @[LZD.scala 39:21]
  wire  _T_1144; // @[LZD.scala 39:30]
  wire  _T_1145; // @[LZD.scala 39:27]
  wire  _T_1146; // @[LZD.scala 39:25]
  wire [1:0] _T_1147; // @[Cat.scala 29:58]
  wire  _T_1148; // @[Shift.scala 12:21]
  wire  _T_1149; // @[Shift.scala 12:21]
  wire  _T_1150; // @[LZD.scala 49:16]
  wire  _T_1151; // @[LZD.scala 49:27]
  wire  _T_1152; // @[LZD.scala 49:25]
  wire  _T_1153; // @[LZD.scala 49:47]
  wire  _T_1154; // @[LZD.scala 49:59]
  wire  _T_1155; // @[LZD.scala 49:35]
  wire [2:0] _T_1157; // @[Cat.scala 29:58]
  wire [3:0] _T_1158; // @[LZD.scala 44:32]
  wire [1:0] _T_1159; // @[LZD.scala 43:32]
  wire  _T_1160; // @[LZD.scala 39:14]
  wire  _T_1161; // @[LZD.scala 39:21]
  wire  _T_1162; // @[LZD.scala 39:30]
  wire  _T_1163; // @[LZD.scala 39:27]
  wire  _T_1164; // @[LZD.scala 39:25]
  wire [1:0] _T_1165; // @[Cat.scala 29:58]
  wire [1:0] _T_1166; // @[LZD.scala 44:32]
  wire  _T_1167; // @[LZD.scala 39:14]
  wire  _T_1168; // @[LZD.scala 39:21]
  wire  _T_1169; // @[LZD.scala 39:30]
  wire  _T_1170; // @[LZD.scala 39:27]
  wire  _T_1171; // @[LZD.scala 39:25]
  wire [1:0] _T_1172; // @[Cat.scala 29:58]
  wire  _T_1173; // @[Shift.scala 12:21]
  wire  _T_1174; // @[Shift.scala 12:21]
  wire  _T_1175; // @[LZD.scala 49:16]
  wire  _T_1176; // @[LZD.scala 49:27]
  wire  _T_1177; // @[LZD.scala 49:25]
  wire  _T_1178; // @[LZD.scala 49:47]
  wire  _T_1179; // @[LZD.scala 49:59]
  wire  _T_1180; // @[LZD.scala 49:35]
  wire [2:0] _T_1182; // @[Cat.scala 29:58]
  wire  _T_1183; // @[Shift.scala 12:21]
  wire  _T_1184; // @[Shift.scala 12:21]
  wire  _T_1185; // @[LZD.scala 49:16]
  wire  _T_1186; // @[LZD.scala 49:27]
  wire  _T_1187; // @[LZD.scala 49:25]
  wire [1:0] _T_1188; // @[LZD.scala 49:47]
  wire [1:0] _T_1189; // @[LZD.scala 49:59]
  wire [1:0] _T_1190; // @[LZD.scala 49:35]
  wire [3:0] _T_1192; // @[Cat.scala 29:58]
  wire  _T_1193; // @[Shift.scala 12:21]
  wire  _T_1194; // @[Shift.scala 12:21]
  wire  _T_1195; // @[LZD.scala 49:16]
  wire  _T_1196; // @[LZD.scala 49:27]
  wire  _T_1197; // @[LZD.scala 49:25]
  wire [2:0] _T_1198; // @[LZD.scala 49:47]
  wire [2:0] _T_1199; // @[LZD.scala 49:59]
  wire [2:0] _T_1200; // @[LZD.scala 49:35]
  wire [4:0] _T_1202; // @[Cat.scala 29:58]
  wire [15:0] _T_1203; // @[LZD.scala 44:32]
  wire [7:0] _T_1204; // @[LZD.scala 43:32]
  wire [3:0] _T_1205; // @[LZD.scala 43:32]
  wire [1:0] _T_1206; // @[LZD.scala 43:32]
  wire  _T_1207; // @[LZD.scala 39:14]
  wire  _T_1208; // @[LZD.scala 39:21]
  wire  _T_1209; // @[LZD.scala 39:30]
  wire  _T_1210; // @[LZD.scala 39:27]
  wire  _T_1211; // @[LZD.scala 39:25]
  wire [1:0] _T_1212; // @[Cat.scala 29:58]
  wire [1:0] _T_1213; // @[LZD.scala 44:32]
  wire  _T_1214; // @[LZD.scala 39:14]
  wire  _T_1215; // @[LZD.scala 39:21]
  wire  _T_1216; // @[LZD.scala 39:30]
  wire  _T_1217; // @[LZD.scala 39:27]
  wire  _T_1218; // @[LZD.scala 39:25]
  wire [1:0] _T_1219; // @[Cat.scala 29:58]
  wire  _T_1220; // @[Shift.scala 12:21]
  wire  _T_1221; // @[Shift.scala 12:21]
  wire  _T_1222; // @[LZD.scala 49:16]
  wire  _T_1223; // @[LZD.scala 49:27]
  wire  _T_1224; // @[LZD.scala 49:25]
  wire  _T_1225; // @[LZD.scala 49:47]
  wire  _T_1226; // @[LZD.scala 49:59]
  wire  _T_1227; // @[LZD.scala 49:35]
  wire [2:0] _T_1229; // @[Cat.scala 29:58]
  wire [3:0] _T_1230; // @[LZD.scala 44:32]
  wire [1:0] _T_1231; // @[LZD.scala 43:32]
  wire  _T_1232; // @[LZD.scala 39:14]
  wire  _T_1233; // @[LZD.scala 39:21]
  wire  _T_1234; // @[LZD.scala 39:30]
  wire  _T_1235; // @[LZD.scala 39:27]
  wire  _T_1236; // @[LZD.scala 39:25]
  wire [1:0] _T_1237; // @[Cat.scala 29:58]
  wire [1:0] _T_1238; // @[LZD.scala 44:32]
  wire  _T_1239; // @[LZD.scala 39:14]
  wire  _T_1240; // @[LZD.scala 39:21]
  wire  _T_1241; // @[LZD.scala 39:30]
  wire  _T_1242; // @[LZD.scala 39:27]
  wire  _T_1243; // @[LZD.scala 39:25]
  wire [1:0] _T_1244; // @[Cat.scala 29:58]
  wire  _T_1245; // @[Shift.scala 12:21]
  wire  _T_1246; // @[Shift.scala 12:21]
  wire  _T_1247; // @[LZD.scala 49:16]
  wire  _T_1248; // @[LZD.scala 49:27]
  wire  _T_1249; // @[LZD.scala 49:25]
  wire  _T_1250; // @[LZD.scala 49:47]
  wire  _T_1251; // @[LZD.scala 49:59]
  wire  _T_1252; // @[LZD.scala 49:35]
  wire [2:0] _T_1254; // @[Cat.scala 29:58]
  wire  _T_1255; // @[Shift.scala 12:21]
  wire  _T_1256; // @[Shift.scala 12:21]
  wire  _T_1257; // @[LZD.scala 49:16]
  wire  _T_1258; // @[LZD.scala 49:27]
  wire  _T_1259; // @[LZD.scala 49:25]
  wire [1:0] _T_1260; // @[LZD.scala 49:47]
  wire [1:0] _T_1261; // @[LZD.scala 49:59]
  wire [1:0] _T_1262; // @[LZD.scala 49:35]
  wire [3:0] _T_1264; // @[Cat.scala 29:58]
  wire [7:0] _T_1265; // @[LZD.scala 44:32]
  wire [3:0] _T_1266; // @[LZD.scala 43:32]
  wire [1:0] _T_1267; // @[LZD.scala 43:32]
  wire  _T_1268; // @[LZD.scala 39:14]
  wire  _T_1269; // @[LZD.scala 39:21]
  wire  _T_1270; // @[LZD.scala 39:30]
  wire  _T_1271; // @[LZD.scala 39:27]
  wire  _T_1272; // @[LZD.scala 39:25]
  wire [1:0] _T_1273; // @[Cat.scala 29:58]
  wire [1:0] _T_1274; // @[LZD.scala 44:32]
  wire  _T_1275; // @[LZD.scala 39:14]
  wire  _T_1276; // @[LZD.scala 39:21]
  wire  _T_1277; // @[LZD.scala 39:30]
  wire  _T_1278; // @[LZD.scala 39:27]
  wire  _T_1279; // @[LZD.scala 39:25]
  wire [1:0] _T_1280; // @[Cat.scala 29:58]
  wire  _T_1281; // @[Shift.scala 12:21]
  wire  _T_1282; // @[Shift.scala 12:21]
  wire  _T_1283; // @[LZD.scala 49:16]
  wire  _T_1284; // @[LZD.scala 49:27]
  wire  _T_1285; // @[LZD.scala 49:25]
  wire  _T_1286; // @[LZD.scala 49:47]
  wire  _T_1287; // @[LZD.scala 49:59]
  wire  _T_1288; // @[LZD.scala 49:35]
  wire [2:0] _T_1290; // @[Cat.scala 29:58]
  wire [3:0] _T_1291; // @[LZD.scala 44:32]
  wire [1:0] _T_1292; // @[LZD.scala 43:32]
  wire  _T_1293; // @[LZD.scala 39:14]
  wire  _T_1294; // @[LZD.scala 39:21]
  wire  _T_1295; // @[LZD.scala 39:30]
  wire  _T_1296; // @[LZD.scala 39:27]
  wire  _T_1297; // @[LZD.scala 39:25]
  wire [1:0] _T_1298; // @[Cat.scala 29:58]
  wire [1:0] _T_1299; // @[LZD.scala 44:32]
  wire  _T_1300; // @[LZD.scala 39:14]
  wire  _T_1301; // @[LZD.scala 39:21]
  wire  _T_1302; // @[LZD.scala 39:30]
  wire  _T_1303; // @[LZD.scala 39:27]
  wire  _T_1304; // @[LZD.scala 39:25]
  wire [1:0] _T_1305; // @[Cat.scala 29:58]
  wire  _T_1306; // @[Shift.scala 12:21]
  wire  _T_1307; // @[Shift.scala 12:21]
  wire  _T_1308; // @[LZD.scala 49:16]
  wire  _T_1309; // @[LZD.scala 49:27]
  wire  _T_1310; // @[LZD.scala 49:25]
  wire  _T_1311; // @[LZD.scala 49:47]
  wire  _T_1312; // @[LZD.scala 49:59]
  wire  _T_1313; // @[LZD.scala 49:35]
  wire [2:0] _T_1315; // @[Cat.scala 29:58]
  wire  _T_1316; // @[Shift.scala 12:21]
  wire  _T_1317; // @[Shift.scala 12:21]
  wire  _T_1318; // @[LZD.scala 49:16]
  wire  _T_1319; // @[LZD.scala 49:27]
  wire  _T_1320; // @[LZD.scala 49:25]
  wire [1:0] _T_1321; // @[LZD.scala 49:47]
  wire [1:0] _T_1322; // @[LZD.scala 49:59]
  wire [1:0] _T_1323; // @[LZD.scala 49:35]
  wire [3:0] _T_1325; // @[Cat.scala 29:58]
  wire  _T_1326; // @[Shift.scala 12:21]
  wire  _T_1327; // @[Shift.scala 12:21]
  wire  _T_1328; // @[LZD.scala 49:16]
  wire  _T_1329; // @[LZD.scala 49:27]
  wire  _T_1330; // @[LZD.scala 49:25]
  wire [2:0] _T_1331; // @[LZD.scala 49:47]
  wire [2:0] _T_1332; // @[LZD.scala 49:59]
  wire [2:0] _T_1333; // @[LZD.scala 49:35]
  wire [4:0] _T_1335; // @[Cat.scala 29:58]
  wire  _T_1336; // @[Shift.scala 12:21]
  wire  _T_1337; // @[Shift.scala 12:21]
  wire  _T_1338; // @[LZD.scala 49:16]
  wire  _T_1339; // @[LZD.scala 49:27]
  wire  _T_1340; // @[LZD.scala 49:25]
  wire [3:0] _T_1341; // @[LZD.scala 49:47]
  wire [3:0] _T_1342; // @[LZD.scala 49:59]
  wire [3:0] _T_1343; // @[LZD.scala 49:35]
  wire [5:0] _T_1345; // @[Cat.scala 29:58]
  wire [26:0] _T_1346; // @[LZD.scala 44:32]
  wire [15:0] _T_1347; // @[LZD.scala 43:32]
  wire [7:0] _T_1348; // @[LZD.scala 43:32]
  wire [3:0] _T_1349; // @[LZD.scala 43:32]
  wire [1:0] _T_1350; // @[LZD.scala 43:32]
  wire  _T_1351; // @[LZD.scala 39:14]
  wire  _T_1352; // @[LZD.scala 39:21]
  wire  _T_1353; // @[LZD.scala 39:30]
  wire  _T_1354; // @[LZD.scala 39:27]
  wire  _T_1355; // @[LZD.scala 39:25]
  wire [1:0] _T_1356; // @[Cat.scala 29:58]
  wire [1:0] _T_1357; // @[LZD.scala 44:32]
  wire  _T_1358; // @[LZD.scala 39:14]
  wire  _T_1359; // @[LZD.scala 39:21]
  wire  _T_1360; // @[LZD.scala 39:30]
  wire  _T_1361; // @[LZD.scala 39:27]
  wire  _T_1362; // @[LZD.scala 39:25]
  wire [1:0] _T_1363; // @[Cat.scala 29:58]
  wire  _T_1364; // @[Shift.scala 12:21]
  wire  _T_1365; // @[Shift.scala 12:21]
  wire  _T_1366; // @[LZD.scala 49:16]
  wire  _T_1367; // @[LZD.scala 49:27]
  wire  _T_1368; // @[LZD.scala 49:25]
  wire  _T_1369; // @[LZD.scala 49:47]
  wire  _T_1370; // @[LZD.scala 49:59]
  wire  _T_1371; // @[LZD.scala 49:35]
  wire [2:0] _T_1373; // @[Cat.scala 29:58]
  wire [3:0] _T_1374; // @[LZD.scala 44:32]
  wire [1:0] _T_1375; // @[LZD.scala 43:32]
  wire  _T_1376; // @[LZD.scala 39:14]
  wire  _T_1377; // @[LZD.scala 39:21]
  wire  _T_1378; // @[LZD.scala 39:30]
  wire  _T_1379; // @[LZD.scala 39:27]
  wire  _T_1380; // @[LZD.scala 39:25]
  wire [1:0] _T_1381; // @[Cat.scala 29:58]
  wire [1:0] _T_1382; // @[LZD.scala 44:32]
  wire  _T_1383; // @[LZD.scala 39:14]
  wire  _T_1384; // @[LZD.scala 39:21]
  wire  _T_1385; // @[LZD.scala 39:30]
  wire  _T_1386; // @[LZD.scala 39:27]
  wire  _T_1387; // @[LZD.scala 39:25]
  wire [1:0] _T_1388; // @[Cat.scala 29:58]
  wire  _T_1389; // @[Shift.scala 12:21]
  wire  _T_1390; // @[Shift.scala 12:21]
  wire  _T_1391; // @[LZD.scala 49:16]
  wire  _T_1392; // @[LZD.scala 49:27]
  wire  _T_1393; // @[LZD.scala 49:25]
  wire  _T_1394; // @[LZD.scala 49:47]
  wire  _T_1395; // @[LZD.scala 49:59]
  wire  _T_1396; // @[LZD.scala 49:35]
  wire [2:0] _T_1398; // @[Cat.scala 29:58]
  wire  _T_1399; // @[Shift.scala 12:21]
  wire  _T_1400; // @[Shift.scala 12:21]
  wire  _T_1401; // @[LZD.scala 49:16]
  wire  _T_1402; // @[LZD.scala 49:27]
  wire  _T_1403; // @[LZD.scala 49:25]
  wire [1:0] _T_1404; // @[LZD.scala 49:47]
  wire [1:0] _T_1405; // @[LZD.scala 49:59]
  wire [1:0] _T_1406; // @[LZD.scala 49:35]
  wire [3:0] _T_1408; // @[Cat.scala 29:58]
  wire [7:0] _T_1409; // @[LZD.scala 44:32]
  wire [3:0] _T_1410; // @[LZD.scala 43:32]
  wire [1:0] _T_1411; // @[LZD.scala 43:32]
  wire  _T_1412; // @[LZD.scala 39:14]
  wire  _T_1413; // @[LZD.scala 39:21]
  wire  _T_1414; // @[LZD.scala 39:30]
  wire  _T_1415; // @[LZD.scala 39:27]
  wire  _T_1416; // @[LZD.scala 39:25]
  wire [1:0] _T_1417; // @[Cat.scala 29:58]
  wire [1:0] _T_1418; // @[LZD.scala 44:32]
  wire  _T_1419; // @[LZD.scala 39:14]
  wire  _T_1420; // @[LZD.scala 39:21]
  wire  _T_1421; // @[LZD.scala 39:30]
  wire  _T_1422; // @[LZD.scala 39:27]
  wire  _T_1423; // @[LZD.scala 39:25]
  wire [1:0] _T_1424; // @[Cat.scala 29:58]
  wire  _T_1425; // @[Shift.scala 12:21]
  wire  _T_1426; // @[Shift.scala 12:21]
  wire  _T_1427; // @[LZD.scala 49:16]
  wire  _T_1428; // @[LZD.scala 49:27]
  wire  _T_1429; // @[LZD.scala 49:25]
  wire  _T_1430; // @[LZD.scala 49:47]
  wire  _T_1431; // @[LZD.scala 49:59]
  wire  _T_1432; // @[LZD.scala 49:35]
  wire [2:0] _T_1434; // @[Cat.scala 29:58]
  wire [3:0] _T_1435; // @[LZD.scala 44:32]
  wire [1:0] _T_1436; // @[LZD.scala 43:32]
  wire  _T_1437; // @[LZD.scala 39:14]
  wire  _T_1438; // @[LZD.scala 39:21]
  wire  _T_1439; // @[LZD.scala 39:30]
  wire  _T_1440; // @[LZD.scala 39:27]
  wire  _T_1441; // @[LZD.scala 39:25]
  wire [1:0] _T_1442; // @[Cat.scala 29:58]
  wire [1:0] _T_1443; // @[LZD.scala 44:32]
  wire  _T_1444; // @[LZD.scala 39:14]
  wire  _T_1445; // @[LZD.scala 39:21]
  wire  _T_1446; // @[LZD.scala 39:30]
  wire  _T_1447; // @[LZD.scala 39:27]
  wire  _T_1448; // @[LZD.scala 39:25]
  wire [1:0] _T_1449; // @[Cat.scala 29:58]
  wire  _T_1450; // @[Shift.scala 12:21]
  wire  _T_1451; // @[Shift.scala 12:21]
  wire  _T_1452; // @[LZD.scala 49:16]
  wire  _T_1453; // @[LZD.scala 49:27]
  wire  _T_1454; // @[LZD.scala 49:25]
  wire  _T_1455; // @[LZD.scala 49:47]
  wire  _T_1456; // @[LZD.scala 49:59]
  wire  _T_1457; // @[LZD.scala 49:35]
  wire [2:0] _T_1459; // @[Cat.scala 29:58]
  wire  _T_1460; // @[Shift.scala 12:21]
  wire  _T_1461; // @[Shift.scala 12:21]
  wire  _T_1462; // @[LZD.scala 49:16]
  wire  _T_1463; // @[LZD.scala 49:27]
  wire  _T_1464; // @[LZD.scala 49:25]
  wire [1:0] _T_1465; // @[LZD.scala 49:47]
  wire [1:0] _T_1466; // @[LZD.scala 49:59]
  wire [1:0] _T_1467; // @[LZD.scala 49:35]
  wire [3:0] _T_1469; // @[Cat.scala 29:58]
  wire  _T_1470; // @[Shift.scala 12:21]
  wire  _T_1471; // @[Shift.scala 12:21]
  wire  _T_1472; // @[LZD.scala 49:16]
  wire  _T_1473; // @[LZD.scala 49:27]
  wire  _T_1474; // @[LZD.scala 49:25]
  wire [2:0] _T_1475; // @[LZD.scala 49:47]
  wire [2:0] _T_1476; // @[LZD.scala 49:59]
  wire [2:0] _T_1477; // @[LZD.scala 49:35]
  wire [4:0] _T_1479; // @[Cat.scala 29:58]
  wire [10:0] _T_1480; // @[LZD.scala 44:32]
  wire [7:0] _T_1481; // @[LZD.scala 43:32]
  wire [3:0] _T_1482; // @[LZD.scala 43:32]
  wire [1:0] _T_1483; // @[LZD.scala 43:32]
  wire  _T_1484; // @[LZD.scala 39:14]
  wire  _T_1485; // @[LZD.scala 39:21]
  wire  _T_1486; // @[LZD.scala 39:30]
  wire  _T_1487; // @[LZD.scala 39:27]
  wire  _T_1488; // @[LZD.scala 39:25]
  wire [1:0] _T_1489; // @[Cat.scala 29:58]
  wire [1:0] _T_1490; // @[LZD.scala 44:32]
  wire  _T_1491; // @[LZD.scala 39:14]
  wire  _T_1492; // @[LZD.scala 39:21]
  wire  _T_1493; // @[LZD.scala 39:30]
  wire  _T_1494; // @[LZD.scala 39:27]
  wire  _T_1495; // @[LZD.scala 39:25]
  wire [1:0] _T_1496; // @[Cat.scala 29:58]
  wire  _T_1497; // @[Shift.scala 12:21]
  wire  _T_1498; // @[Shift.scala 12:21]
  wire  _T_1499; // @[LZD.scala 49:16]
  wire  _T_1500; // @[LZD.scala 49:27]
  wire  _T_1501; // @[LZD.scala 49:25]
  wire  _T_1502; // @[LZD.scala 49:47]
  wire  _T_1503; // @[LZD.scala 49:59]
  wire  _T_1504; // @[LZD.scala 49:35]
  wire [2:0] _T_1506; // @[Cat.scala 29:58]
  wire [3:0] _T_1507; // @[LZD.scala 44:32]
  wire [1:0] _T_1508; // @[LZD.scala 43:32]
  wire  _T_1509; // @[LZD.scala 39:14]
  wire  _T_1510; // @[LZD.scala 39:21]
  wire  _T_1511; // @[LZD.scala 39:30]
  wire  _T_1512; // @[LZD.scala 39:27]
  wire  _T_1513; // @[LZD.scala 39:25]
  wire [1:0] _T_1514; // @[Cat.scala 29:58]
  wire [1:0] _T_1515; // @[LZD.scala 44:32]
  wire  _T_1516; // @[LZD.scala 39:14]
  wire  _T_1517; // @[LZD.scala 39:21]
  wire  _T_1518; // @[LZD.scala 39:30]
  wire  _T_1519; // @[LZD.scala 39:27]
  wire  _T_1520; // @[LZD.scala 39:25]
  wire [1:0] _T_1521; // @[Cat.scala 29:58]
  wire  _T_1522; // @[Shift.scala 12:21]
  wire  _T_1523; // @[Shift.scala 12:21]
  wire  _T_1524; // @[LZD.scala 49:16]
  wire  _T_1525; // @[LZD.scala 49:27]
  wire  _T_1526; // @[LZD.scala 49:25]
  wire  _T_1527; // @[LZD.scala 49:47]
  wire  _T_1528; // @[LZD.scala 49:59]
  wire  _T_1529; // @[LZD.scala 49:35]
  wire [2:0] _T_1531; // @[Cat.scala 29:58]
  wire  _T_1532; // @[Shift.scala 12:21]
  wire  _T_1533; // @[Shift.scala 12:21]
  wire  _T_1534; // @[LZD.scala 49:16]
  wire  _T_1535; // @[LZD.scala 49:27]
  wire  _T_1536; // @[LZD.scala 49:25]
  wire [1:0] _T_1537; // @[LZD.scala 49:47]
  wire [1:0] _T_1538; // @[LZD.scala 49:59]
  wire [1:0] _T_1539; // @[LZD.scala 49:35]
  wire [3:0] _T_1541; // @[Cat.scala 29:58]
  wire [2:0] _T_1542; // @[LZD.scala 44:32]
  wire [1:0] _T_1543; // @[LZD.scala 43:32]
  wire  _T_1544; // @[LZD.scala 39:14]
  wire  _T_1545; // @[LZD.scala 39:21]
  wire  _T_1546; // @[LZD.scala 39:30]
  wire  _T_1547; // @[LZD.scala 39:27]
  wire  _T_1548; // @[LZD.scala 39:25]
  wire [1:0] _T_1549; // @[Cat.scala 29:58]
  wire  _T_1550; // @[LZD.scala 44:32]
  wire  _T_1552; // @[Shift.scala 12:21]
  wire  _T_1554; // @[LZD.scala 55:32]
  wire  _T_1555; // @[LZD.scala 55:20]
  wire  _T_1557; // @[Shift.scala 12:21]
  wire [2:0] _T_1559; // @[Cat.scala 29:58]
  wire [2:0] _T_1560; // @[LZD.scala 55:32]
  wire [2:0] _T_1561; // @[LZD.scala 55:20]
  wire [3:0] _T_1562; // @[Cat.scala 29:58]
  wire  _T_1563; // @[Shift.scala 12:21]
  wire [3:0] _T_1565; // @[LZD.scala 55:32]
  wire [3:0] _T_1566; // @[LZD.scala 55:20]
  wire [4:0] _T_1567; // @[Cat.scala 29:58]
  wire  _T_1568; // @[Shift.scala 12:21]
  wire [4:0] _T_1570; // @[LZD.scala 55:32]
  wire [4:0] _T_1571; // @[LZD.scala 55:20]
  wire [5:0] sumLZD; // @[Cat.scala 29:58]
  wire [5:0] shiftValue; // @[PositFMA.scala 126:24]
  wire [57:0] _T_1572; // @[PositFMA.scala 127:38]
  wire  _T_1573; // @[Shift.scala 16:24]
  wire  _T_1575; // @[Shift.scala 12:21]
  wire [25:0] _T_1576; // @[Shift.scala 64:52]
  wire [57:0] _T_1578; // @[Cat.scala 29:58]
  wire [57:0] _T_1579; // @[Shift.scala 64:27]
  wire [4:0] _T_1580; // @[Shift.scala 66:70]
  wire  _T_1581; // @[Shift.scala 12:21]
  wire [41:0] _T_1582; // @[Shift.scala 64:52]
  wire [57:0] _T_1584; // @[Cat.scala 29:58]
  wire [57:0] _T_1585; // @[Shift.scala 64:27]
  wire [3:0] _T_1586; // @[Shift.scala 66:70]
  wire  _T_1587; // @[Shift.scala 12:21]
  wire [49:0] _T_1588; // @[Shift.scala 64:52]
  wire [57:0] _T_1590; // @[Cat.scala 29:58]
  wire [57:0] _T_1591; // @[Shift.scala 64:27]
  wire [2:0] _T_1592; // @[Shift.scala 66:70]
  wire  _T_1593; // @[Shift.scala 12:21]
  wire [53:0] _T_1594; // @[Shift.scala 64:52]
  wire [57:0] _T_1596; // @[Cat.scala 29:58]
  wire [57:0] _T_1597; // @[Shift.scala 64:27]
  wire [1:0] _T_1598; // @[Shift.scala 66:70]
  wire  _T_1599; // @[Shift.scala 12:21]
  wire [55:0] _T_1600; // @[Shift.scala 64:52]
  wire [57:0] _T_1602; // @[Cat.scala 29:58]
  wire [57:0] _T_1603; // @[Shift.scala 64:27]
  wire  _T_1604; // @[Shift.scala 66:70]
  wire [56:0] _T_1606; // @[Shift.scala 64:52]
  wire [57:0] _T_1607; // @[Cat.scala 29:58]
  wire [57:0] _T_1608; // @[Shift.scala 64:27]
  wire [57:0] normalFracTmp; // @[Shift.scala 16:10]
  wire [7:0] _T_1610; // @[PositFMA.scala 130:36]
  wire [7:0] _T_1611; // @[PositFMA.scala 130:36]
  wire [6:0] _T_1612; // @[Cat.scala 29:58]
  wire [6:0] _T_1613; // @[PositFMA.scala 130:61]
  wire [7:0] _GEN_20; // @[PositFMA.scala 130:42]
  wire [7:0] _T_1615; // @[PositFMA.scala 130:42]
  wire [7:0] sumScale; // @[PositFMA.scala 130:42]
  wire [27:0] sumFrac; // @[PositFMA.scala 131:41]
  wire [29:0] grsTmp; // @[PositFMA.scala 134:41]
  wire [1:0] _T_1616; // @[PositFMA.scala 137:40]
  wire [27:0] _T_1617; // @[PositFMA.scala 137:56]
  wire  _T_1618; // @[PositFMA.scala 137:60]
  wire  underflow; // @[PositFMA.scala 144:32]
  wire  overflow; // @[PositFMA.scala 145:32]
  wire  _T_1619; // @[PositFMA.scala 154:32]
  wire  decF_isZero; // @[PositFMA.scala 154:20]
  wire [7:0] _T_1621; // @[Mux.scala 87:16]
  wire [7:0] _T_1622; // @[Mux.scala 87:16]
  wire [6:0] _GEN_21; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  wire [6:0] decF_scale; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  wire  _T_1623; // @[convert.scala 46:61]
  wire  _T_1624; // @[convert.scala 46:52]
  wire  _T_1626; // @[convert.scala 46:42]
  wire [5:0] _T_1627; // @[convert.scala 48:34]
  wire  _T_1628; // @[convert.scala 49:36]
  wire [5:0] _T_1630; // @[convert.scala 50:36]
  wire [5:0] _T_1631; // @[convert.scala 50:36]
  wire [5:0] _T_1632; // @[convert.scala 50:28]
  wire  _T_1633; // @[convert.scala 51:31]
  wire  _T_1634; // @[convert.scala 52:43]
  wire [33:0] _T_1638; // @[Cat.scala 29:58]
  wire [5:0] _T_1639; // @[Shift.scala 39:17]
  wire  _T_1640; // @[Shift.scala 39:24]
  wire [1:0] _T_1642; // @[Shift.scala 90:30]
  wire [31:0] _T_1643; // @[Shift.scala 90:48]
  wire  _T_1644; // @[Shift.scala 90:57]
  wire [1:0] _GEN_22; // @[Shift.scala 90:39]
  wire [1:0] _T_1645; // @[Shift.scala 90:39]
  wire  _T_1646; // @[Shift.scala 12:21]
  wire  _T_1647; // @[Shift.scala 12:21]
  wire [31:0] _T_1649; // @[Bitwise.scala 71:12]
  wire [33:0] _T_1650; // @[Cat.scala 29:58]
  wire [33:0] _T_1651; // @[Shift.scala 91:22]
  wire [4:0] _T_1652; // @[Shift.scala 92:77]
  wire [17:0] _T_1653; // @[Shift.scala 90:30]
  wire [15:0] _T_1654; // @[Shift.scala 90:48]
  wire  _T_1655; // @[Shift.scala 90:57]
  wire [17:0] _GEN_23; // @[Shift.scala 90:39]
  wire [17:0] _T_1656; // @[Shift.scala 90:39]
  wire  _T_1657; // @[Shift.scala 12:21]
  wire  _T_1658; // @[Shift.scala 12:21]
  wire [15:0] _T_1660; // @[Bitwise.scala 71:12]
  wire [33:0] _T_1661; // @[Cat.scala 29:58]
  wire [33:0] _T_1662; // @[Shift.scala 91:22]
  wire [3:0] _T_1663; // @[Shift.scala 92:77]
  wire [25:0] _T_1664; // @[Shift.scala 90:30]
  wire [7:0] _T_1665; // @[Shift.scala 90:48]
  wire  _T_1666; // @[Shift.scala 90:57]
  wire [25:0] _GEN_24; // @[Shift.scala 90:39]
  wire [25:0] _T_1667; // @[Shift.scala 90:39]
  wire  _T_1668; // @[Shift.scala 12:21]
  wire  _T_1669; // @[Shift.scala 12:21]
  wire [7:0] _T_1671; // @[Bitwise.scala 71:12]
  wire [33:0] _T_1672; // @[Cat.scala 29:58]
  wire [33:0] _T_1673; // @[Shift.scala 91:22]
  wire [2:0] _T_1674; // @[Shift.scala 92:77]
  wire [29:0] _T_1675; // @[Shift.scala 90:30]
  wire [3:0] _T_1676; // @[Shift.scala 90:48]
  wire  _T_1677; // @[Shift.scala 90:57]
  wire [29:0] _GEN_25; // @[Shift.scala 90:39]
  wire [29:0] _T_1678; // @[Shift.scala 90:39]
  wire  _T_1679; // @[Shift.scala 12:21]
  wire  _T_1680; // @[Shift.scala 12:21]
  wire [3:0] _T_1682; // @[Bitwise.scala 71:12]
  wire [33:0] _T_1683; // @[Cat.scala 29:58]
  wire [33:0] _T_1684; // @[Shift.scala 91:22]
  wire [1:0] _T_1685; // @[Shift.scala 92:77]
  wire [31:0] _T_1686; // @[Shift.scala 90:30]
  wire [1:0] _T_1687; // @[Shift.scala 90:48]
  wire  _T_1688; // @[Shift.scala 90:57]
  wire [31:0] _GEN_26; // @[Shift.scala 90:39]
  wire [31:0] _T_1689; // @[Shift.scala 90:39]
  wire  _T_1690; // @[Shift.scala 12:21]
  wire  _T_1691; // @[Shift.scala 12:21]
  wire [1:0] _T_1693; // @[Bitwise.scala 71:12]
  wire [33:0] _T_1694; // @[Cat.scala 29:58]
  wire [33:0] _T_1695; // @[Shift.scala 91:22]
  wire  _T_1696; // @[Shift.scala 92:77]
  wire [32:0] _T_1697; // @[Shift.scala 90:30]
  wire  _T_1698; // @[Shift.scala 90:48]
  wire [32:0] _GEN_27; // @[Shift.scala 90:39]
  wire [32:0] _T_1700; // @[Shift.scala 90:39]
  wire  _T_1702; // @[Shift.scala 12:21]
  wire [33:0] _T_1703; // @[Cat.scala 29:58]
  wire [33:0] _T_1704; // @[Shift.scala 91:22]
  wire [33:0] _T_1707; // @[Bitwise.scala 71:12]
  wire [33:0] _T_1708; // @[Shift.scala 39:10]
  wire  _T_1709; // @[convert.scala 55:31]
  wire  _T_1710; // @[convert.scala 56:31]
  wire  _T_1711; // @[convert.scala 57:31]
  wire  _T_1712; // @[convert.scala 58:31]
  wire [30:0] _T_1713; // @[convert.scala 59:69]
  wire  _T_1714; // @[convert.scala 59:81]
  wire  _T_1715; // @[convert.scala 59:50]
  wire  _T_1717; // @[convert.scala 60:81]
  wire  _T_1718; // @[convert.scala 61:44]
  wire  _T_1719; // @[convert.scala 61:52]
  wire  _T_1720; // @[convert.scala 61:36]
  wire  _T_1721; // @[convert.scala 62:63]
  wire  _T_1722; // @[convert.scala 62:103]
  wire  _T_1723; // @[convert.scala 62:60]
  wire [30:0] _GEN_28; // @[convert.scala 63:56]
  wire [30:0] _T_1726; // @[convert.scala 63:56]
  wire [31:0] _T_1727; // @[Cat.scala 29:58]
  reg  _T_1731; // @[Valid.scala 117:22]
  reg [31:0] _RAND_8;
  reg [31:0] _T_1735; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  assign _T = io_fmaOp[1]; // @[PositFMA.scala 47:36]
  assign _T_2 = _T ? 32'hffffffff : 32'h0; // @[Bitwise.scala 71:12]
  assign _T_3 = _T_2 ^ io_A; // @[PositFMA.scala 47:41]
  assign _GEN_10 = {{31'd0}, _T}; // @[PositFMA.scala 47:49]
  assign realA = _T_3 + _GEN_10; // @[PositFMA.scala 47:49]
  assign _T_6 = io_fmaOp[0]; // @[PositFMA.scala 48:36]
  assign _T_8 = _T_6 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 71:12]
  assign _T_9 = _T_8 ^ io_C; // @[PositFMA.scala 48:41]
  assign _GEN_11 = {{31'd0}, _T_6}; // @[PositFMA.scala 48:49]
  assign realC = _T_9 + _GEN_11; // @[PositFMA.scala 48:49]
  assign _T_13 = realA[31]; // @[convert.scala 18:24]
  assign _T_14 = realA[30]; // @[convert.scala 18:40]
  assign _T_15 = _T_13 ^ _T_14; // @[convert.scala 18:36]
  assign _T_16 = realA[30:1]; // @[convert.scala 19:24]
  assign _T_17 = realA[29:0]; // @[convert.scala 19:43]
  assign _T_18 = _T_16 ^ _T_17; // @[convert.scala 19:39]
  assign _T_19 = _T_18[29:14]; // @[LZD.scala 43:32]
  assign _T_20 = _T_19[15:8]; // @[LZD.scala 43:32]
  assign _T_21 = _T_20[7:4]; // @[LZD.scala 43:32]
  assign _T_22 = _T_21[3:2]; // @[LZD.scala 43:32]
  assign _T_23 = _T_22 != 2'h0; // @[LZD.scala 39:14]
  assign _T_24 = _T_22[1]; // @[LZD.scala 39:21]
  assign _T_25 = _T_22[0]; // @[LZD.scala 39:30]
  assign _T_26 = ~ _T_25; // @[LZD.scala 39:27]
  assign _T_27 = _T_24 | _T_26; // @[LZD.scala 39:25]
  assign _T_28 = {_T_23,_T_27}; // @[Cat.scala 29:58]
  assign _T_29 = _T_21[1:0]; // @[LZD.scala 44:32]
  assign _T_30 = _T_29 != 2'h0; // @[LZD.scala 39:14]
  assign _T_31 = _T_29[1]; // @[LZD.scala 39:21]
  assign _T_32 = _T_29[0]; // @[LZD.scala 39:30]
  assign _T_33 = ~ _T_32; // @[LZD.scala 39:27]
  assign _T_34 = _T_31 | _T_33; // @[LZD.scala 39:25]
  assign _T_35 = {_T_30,_T_34}; // @[Cat.scala 29:58]
  assign _T_36 = _T_28[1]; // @[Shift.scala 12:21]
  assign _T_37 = _T_35[1]; // @[Shift.scala 12:21]
  assign _T_38 = _T_36 | _T_37; // @[LZD.scala 49:16]
  assign _T_39 = ~ _T_37; // @[LZD.scala 49:27]
  assign _T_40 = _T_36 | _T_39; // @[LZD.scala 49:25]
  assign _T_41 = _T_28[0:0]; // @[LZD.scala 49:47]
  assign _T_42 = _T_35[0:0]; // @[LZD.scala 49:59]
  assign _T_43 = _T_36 ? _T_41 : _T_42; // @[LZD.scala 49:35]
  assign _T_45 = {_T_38,_T_40,_T_43}; // @[Cat.scala 29:58]
  assign _T_46 = _T_20[3:0]; // @[LZD.scala 44:32]
  assign _T_47 = _T_46[3:2]; // @[LZD.scala 43:32]
  assign _T_48 = _T_47 != 2'h0; // @[LZD.scala 39:14]
  assign _T_49 = _T_47[1]; // @[LZD.scala 39:21]
  assign _T_50 = _T_47[0]; // @[LZD.scala 39:30]
  assign _T_51 = ~ _T_50; // @[LZD.scala 39:27]
  assign _T_52 = _T_49 | _T_51; // @[LZD.scala 39:25]
  assign _T_53 = {_T_48,_T_52}; // @[Cat.scala 29:58]
  assign _T_54 = _T_46[1:0]; // @[LZD.scala 44:32]
  assign _T_55 = _T_54 != 2'h0; // @[LZD.scala 39:14]
  assign _T_56 = _T_54[1]; // @[LZD.scala 39:21]
  assign _T_57 = _T_54[0]; // @[LZD.scala 39:30]
  assign _T_58 = ~ _T_57; // @[LZD.scala 39:27]
  assign _T_59 = _T_56 | _T_58; // @[LZD.scala 39:25]
  assign _T_60 = {_T_55,_T_59}; // @[Cat.scala 29:58]
  assign _T_61 = _T_53[1]; // @[Shift.scala 12:21]
  assign _T_62 = _T_60[1]; // @[Shift.scala 12:21]
  assign _T_63 = _T_61 | _T_62; // @[LZD.scala 49:16]
  assign _T_64 = ~ _T_62; // @[LZD.scala 49:27]
  assign _T_65 = _T_61 | _T_64; // @[LZD.scala 49:25]
  assign _T_66 = _T_53[0:0]; // @[LZD.scala 49:47]
  assign _T_67 = _T_60[0:0]; // @[LZD.scala 49:59]
  assign _T_68 = _T_61 ? _T_66 : _T_67; // @[LZD.scala 49:35]
  assign _T_70 = {_T_63,_T_65,_T_68}; // @[Cat.scala 29:58]
  assign _T_71 = _T_45[2]; // @[Shift.scala 12:21]
  assign _T_72 = _T_70[2]; // @[Shift.scala 12:21]
  assign _T_73 = _T_71 | _T_72; // @[LZD.scala 49:16]
  assign _T_74 = ~ _T_72; // @[LZD.scala 49:27]
  assign _T_75 = _T_71 | _T_74; // @[LZD.scala 49:25]
  assign _T_76 = _T_45[1:0]; // @[LZD.scala 49:47]
  assign _T_77 = _T_70[1:0]; // @[LZD.scala 49:59]
  assign _T_78 = _T_71 ? _T_76 : _T_77; // @[LZD.scala 49:35]
  assign _T_80 = {_T_73,_T_75,_T_78}; // @[Cat.scala 29:58]
  assign _T_81 = _T_19[7:0]; // @[LZD.scala 44:32]
  assign _T_82 = _T_81[7:4]; // @[LZD.scala 43:32]
  assign _T_83 = _T_82[3:2]; // @[LZD.scala 43:32]
  assign _T_84 = _T_83 != 2'h0; // @[LZD.scala 39:14]
  assign _T_85 = _T_83[1]; // @[LZD.scala 39:21]
  assign _T_86 = _T_83[0]; // @[LZD.scala 39:30]
  assign _T_87 = ~ _T_86; // @[LZD.scala 39:27]
  assign _T_88 = _T_85 | _T_87; // @[LZD.scala 39:25]
  assign _T_89 = {_T_84,_T_88}; // @[Cat.scala 29:58]
  assign _T_90 = _T_82[1:0]; // @[LZD.scala 44:32]
  assign _T_91 = _T_90 != 2'h0; // @[LZD.scala 39:14]
  assign _T_92 = _T_90[1]; // @[LZD.scala 39:21]
  assign _T_93 = _T_90[0]; // @[LZD.scala 39:30]
  assign _T_94 = ~ _T_93; // @[LZD.scala 39:27]
  assign _T_95 = _T_92 | _T_94; // @[LZD.scala 39:25]
  assign _T_96 = {_T_91,_T_95}; // @[Cat.scala 29:58]
  assign _T_97 = _T_89[1]; // @[Shift.scala 12:21]
  assign _T_98 = _T_96[1]; // @[Shift.scala 12:21]
  assign _T_99 = _T_97 | _T_98; // @[LZD.scala 49:16]
  assign _T_100 = ~ _T_98; // @[LZD.scala 49:27]
  assign _T_101 = _T_97 | _T_100; // @[LZD.scala 49:25]
  assign _T_102 = _T_89[0:0]; // @[LZD.scala 49:47]
  assign _T_103 = _T_96[0:0]; // @[LZD.scala 49:59]
  assign _T_104 = _T_97 ? _T_102 : _T_103; // @[LZD.scala 49:35]
  assign _T_106 = {_T_99,_T_101,_T_104}; // @[Cat.scala 29:58]
  assign _T_107 = _T_81[3:0]; // @[LZD.scala 44:32]
  assign _T_108 = _T_107[3:2]; // @[LZD.scala 43:32]
  assign _T_109 = _T_108 != 2'h0; // @[LZD.scala 39:14]
  assign _T_110 = _T_108[1]; // @[LZD.scala 39:21]
  assign _T_111 = _T_108[0]; // @[LZD.scala 39:30]
  assign _T_112 = ~ _T_111; // @[LZD.scala 39:27]
  assign _T_113 = _T_110 | _T_112; // @[LZD.scala 39:25]
  assign _T_114 = {_T_109,_T_113}; // @[Cat.scala 29:58]
  assign _T_115 = _T_107[1:0]; // @[LZD.scala 44:32]
  assign _T_116 = _T_115 != 2'h0; // @[LZD.scala 39:14]
  assign _T_117 = _T_115[1]; // @[LZD.scala 39:21]
  assign _T_118 = _T_115[0]; // @[LZD.scala 39:30]
  assign _T_119 = ~ _T_118; // @[LZD.scala 39:27]
  assign _T_120 = _T_117 | _T_119; // @[LZD.scala 39:25]
  assign _T_121 = {_T_116,_T_120}; // @[Cat.scala 29:58]
  assign _T_122 = _T_114[1]; // @[Shift.scala 12:21]
  assign _T_123 = _T_121[1]; // @[Shift.scala 12:21]
  assign _T_124 = _T_122 | _T_123; // @[LZD.scala 49:16]
  assign _T_125 = ~ _T_123; // @[LZD.scala 49:27]
  assign _T_126 = _T_122 | _T_125; // @[LZD.scala 49:25]
  assign _T_127 = _T_114[0:0]; // @[LZD.scala 49:47]
  assign _T_128 = _T_121[0:0]; // @[LZD.scala 49:59]
  assign _T_129 = _T_122 ? _T_127 : _T_128; // @[LZD.scala 49:35]
  assign _T_131 = {_T_124,_T_126,_T_129}; // @[Cat.scala 29:58]
  assign _T_132 = _T_106[2]; // @[Shift.scala 12:21]
  assign _T_133 = _T_131[2]; // @[Shift.scala 12:21]
  assign _T_134 = _T_132 | _T_133; // @[LZD.scala 49:16]
  assign _T_135 = ~ _T_133; // @[LZD.scala 49:27]
  assign _T_136 = _T_132 | _T_135; // @[LZD.scala 49:25]
  assign _T_137 = _T_106[1:0]; // @[LZD.scala 49:47]
  assign _T_138 = _T_131[1:0]; // @[LZD.scala 49:59]
  assign _T_139 = _T_132 ? _T_137 : _T_138; // @[LZD.scala 49:35]
  assign _T_141 = {_T_134,_T_136,_T_139}; // @[Cat.scala 29:58]
  assign _T_142 = _T_80[3]; // @[Shift.scala 12:21]
  assign _T_143 = _T_141[3]; // @[Shift.scala 12:21]
  assign _T_144 = _T_142 | _T_143; // @[LZD.scala 49:16]
  assign _T_145 = ~ _T_143; // @[LZD.scala 49:27]
  assign _T_146 = _T_142 | _T_145; // @[LZD.scala 49:25]
  assign _T_147 = _T_80[2:0]; // @[LZD.scala 49:47]
  assign _T_148 = _T_141[2:0]; // @[LZD.scala 49:59]
  assign _T_149 = _T_142 ? _T_147 : _T_148; // @[LZD.scala 49:35]
  assign _T_151 = {_T_144,_T_146,_T_149}; // @[Cat.scala 29:58]
  assign _T_152 = _T_18[13:0]; // @[LZD.scala 44:32]
  assign _T_153 = _T_152[13:6]; // @[LZD.scala 43:32]
  assign _T_154 = _T_153[7:4]; // @[LZD.scala 43:32]
  assign _T_155 = _T_154[3:2]; // @[LZD.scala 43:32]
  assign _T_156 = _T_155 != 2'h0; // @[LZD.scala 39:14]
  assign _T_157 = _T_155[1]; // @[LZD.scala 39:21]
  assign _T_158 = _T_155[0]; // @[LZD.scala 39:30]
  assign _T_159 = ~ _T_158; // @[LZD.scala 39:27]
  assign _T_160 = _T_157 | _T_159; // @[LZD.scala 39:25]
  assign _T_161 = {_T_156,_T_160}; // @[Cat.scala 29:58]
  assign _T_162 = _T_154[1:0]; // @[LZD.scala 44:32]
  assign _T_163 = _T_162 != 2'h0; // @[LZD.scala 39:14]
  assign _T_164 = _T_162[1]; // @[LZD.scala 39:21]
  assign _T_165 = _T_162[0]; // @[LZD.scala 39:30]
  assign _T_166 = ~ _T_165; // @[LZD.scala 39:27]
  assign _T_167 = _T_164 | _T_166; // @[LZD.scala 39:25]
  assign _T_168 = {_T_163,_T_167}; // @[Cat.scala 29:58]
  assign _T_169 = _T_161[1]; // @[Shift.scala 12:21]
  assign _T_170 = _T_168[1]; // @[Shift.scala 12:21]
  assign _T_171 = _T_169 | _T_170; // @[LZD.scala 49:16]
  assign _T_172 = ~ _T_170; // @[LZD.scala 49:27]
  assign _T_173 = _T_169 | _T_172; // @[LZD.scala 49:25]
  assign _T_174 = _T_161[0:0]; // @[LZD.scala 49:47]
  assign _T_175 = _T_168[0:0]; // @[LZD.scala 49:59]
  assign _T_176 = _T_169 ? _T_174 : _T_175; // @[LZD.scala 49:35]
  assign _T_178 = {_T_171,_T_173,_T_176}; // @[Cat.scala 29:58]
  assign _T_179 = _T_153[3:0]; // @[LZD.scala 44:32]
  assign _T_180 = _T_179[3:2]; // @[LZD.scala 43:32]
  assign _T_181 = _T_180 != 2'h0; // @[LZD.scala 39:14]
  assign _T_182 = _T_180[1]; // @[LZD.scala 39:21]
  assign _T_183 = _T_180[0]; // @[LZD.scala 39:30]
  assign _T_184 = ~ _T_183; // @[LZD.scala 39:27]
  assign _T_185 = _T_182 | _T_184; // @[LZD.scala 39:25]
  assign _T_186 = {_T_181,_T_185}; // @[Cat.scala 29:58]
  assign _T_187 = _T_179[1:0]; // @[LZD.scala 44:32]
  assign _T_188 = _T_187 != 2'h0; // @[LZD.scala 39:14]
  assign _T_189 = _T_187[1]; // @[LZD.scala 39:21]
  assign _T_190 = _T_187[0]; // @[LZD.scala 39:30]
  assign _T_191 = ~ _T_190; // @[LZD.scala 39:27]
  assign _T_192 = _T_189 | _T_191; // @[LZD.scala 39:25]
  assign _T_193 = {_T_188,_T_192}; // @[Cat.scala 29:58]
  assign _T_194 = _T_186[1]; // @[Shift.scala 12:21]
  assign _T_195 = _T_193[1]; // @[Shift.scala 12:21]
  assign _T_196 = _T_194 | _T_195; // @[LZD.scala 49:16]
  assign _T_197 = ~ _T_195; // @[LZD.scala 49:27]
  assign _T_198 = _T_194 | _T_197; // @[LZD.scala 49:25]
  assign _T_199 = _T_186[0:0]; // @[LZD.scala 49:47]
  assign _T_200 = _T_193[0:0]; // @[LZD.scala 49:59]
  assign _T_201 = _T_194 ? _T_199 : _T_200; // @[LZD.scala 49:35]
  assign _T_203 = {_T_196,_T_198,_T_201}; // @[Cat.scala 29:58]
  assign _T_204 = _T_178[2]; // @[Shift.scala 12:21]
  assign _T_205 = _T_203[2]; // @[Shift.scala 12:21]
  assign _T_206 = _T_204 | _T_205; // @[LZD.scala 49:16]
  assign _T_207 = ~ _T_205; // @[LZD.scala 49:27]
  assign _T_208 = _T_204 | _T_207; // @[LZD.scala 49:25]
  assign _T_209 = _T_178[1:0]; // @[LZD.scala 49:47]
  assign _T_210 = _T_203[1:0]; // @[LZD.scala 49:59]
  assign _T_211 = _T_204 ? _T_209 : _T_210; // @[LZD.scala 49:35]
  assign _T_213 = {_T_206,_T_208,_T_211}; // @[Cat.scala 29:58]
  assign _T_214 = _T_152[5:0]; // @[LZD.scala 44:32]
  assign _T_215 = _T_214[5:2]; // @[LZD.scala 43:32]
  assign _T_216 = _T_215[3:2]; // @[LZD.scala 43:32]
  assign _T_217 = _T_216 != 2'h0; // @[LZD.scala 39:14]
  assign _T_218 = _T_216[1]; // @[LZD.scala 39:21]
  assign _T_219 = _T_216[0]; // @[LZD.scala 39:30]
  assign _T_220 = ~ _T_219; // @[LZD.scala 39:27]
  assign _T_221 = _T_218 | _T_220; // @[LZD.scala 39:25]
  assign _T_222 = {_T_217,_T_221}; // @[Cat.scala 29:58]
  assign _T_223 = _T_215[1:0]; // @[LZD.scala 44:32]
  assign _T_224 = _T_223 != 2'h0; // @[LZD.scala 39:14]
  assign _T_225 = _T_223[1]; // @[LZD.scala 39:21]
  assign _T_226 = _T_223[0]; // @[LZD.scala 39:30]
  assign _T_227 = ~ _T_226; // @[LZD.scala 39:27]
  assign _T_228 = _T_225 | _T_227; // @[LZD.scala 39:25]
  assign _T_229 = {_T_224,_T_228}; // @[Cat.scala 29:58]
  assign _T_230 = _T_222[1]; // @[Shift.scala 12:21]
  assign _T_231 = _T_229[1]; // @[Shift.scala 12:21]
  assign _T_232 = _T_230 | _T_231; // @[LZD.scala 49:16]
  assign _T_233 = ~ _T_231; // @[LZD.scala 49:27]
  assign _T_234 = _T_230 | _T_233; // @[LZD.scala 49:25]
  assign _T_235 = _T_222[0:0]; // @[LZD.scala 49:47]
  assign _T_236 = _T_229[0:0]; // @[LZD.scala 49:59]
  assign _T_237 = _T_230 ? _T_235 : _T_236; // @[LZD.scala 49:35]
  assign _T_239 = {_T_232,_T_234,_T_237}; // @[Cat.scala 29:58]
  assign _T_240 = _T_214[1:0]; // @[LZD.scala 44:32]
  assign _T_241 = _T_240 != 2'h0; // @[LZD.scala 39:14]
  assign _T_242 = _T_240[1]; // @[LZD.scala 39:21]
  assign _T_243 = _T_240[0]; // @[LZD.scala 39:30]
  assign _T_244 = ~ _T_243; // @[LZD.scala 39:27]
  assign _T_245 = _T_242 | _T_244; // @[LZD.scala 39:25]
  assign _T_246 = {_T_241,_T_245}; // @[Cat.scala 29:58]
  assign _T_247 = _T_239[2]; // @[Shift.scala 12:21]
  assign _T_249 = _T_239[1:0]; // @[LZD.scala 55:32]
  assign _T_250 = _T_247 ? _T_249 : _T_246; // @[LZD.scala 55:20]
  assign _T_251 = {_T_247,_T_250}; // @[Cat.scala 29:58]
  assign _T_252 = _T_213[3]; // @[Shift.scala 12:21]
  assign _T_254 = _T_213[2:0]; // @[LZD.scala 55:32]
  assign _T_255 = _T_252 ? _T_254 : _T_251; // @[LZD.scala 55:20]
  assign _T_256 = {_T_252,_T_255}; // @[Cat.scala 29:58]
  assign _T_257 = _T_151[4]; // @[Shift.scala 12:21]
  assign _T_259 = _T_151[3:0]; // @[LZD.scala 55:32]
  assign _T_260 = _T_257 ? _T_259 : _T_256; // @[LZD.scala 55:20]
  assign _T_261 = {_T_257,_T_260}; // @[Cat.scala 29:58]
  assign _T_262 = ~ _T_261; // @[convert.scala 21:22]
  assign _T_263 = realA[28:0]; // @[convert.scala 22:36]
  assign _T_264 = _T_262 < 5'h1d; // @[Shift.scala 16:24]
  assign _T_266 = _T_262[4]; // @[Shift.scala 12:21]
  assign _T_267 = _T_263[12:0]; // @[Shift.scala 64:52]
  assign _T_269 = {_T_267,16'h0}; // @[Cat.scala 29:58]
  assign _T_270 = _T_266 ? _T_269 : _T_263; // @[Shift.scala 64:27]
  assign _T_271 = _T_262[3:0]; // @[Shift.scala 66:70]
  assign _T_272 = _T_271[3]; // @[Shift.scala 12:21]
  assign _T_273 = _T_270[20:0]; // @[Shift.scala 64:52]
  assign _T_275 = {_T_273,8'h0}; // @[Cat.scala 29:58]
  assign _T_276 = _T_272 ? _T_275 : _T_270; // @[Shift.scala 64:27]
  assign _T_277 = _T_271[2:0]; // @[Shift.scala 66:70]
  assign _T_278 = _T_277[2]; // @[Shift.scala 12:21]
  assign _T_279 = _T_276[24:0]; // @[Shift.scala 64:52]
  assign _T_281 = {_T_279,4'h0}; // @[Cat.scala 29:58]
  assign _T_282 = _T_278 ? _T_281 : _T_276; // @[Shift.scala 64:27]
  assign _T_283 = _T_277[1:0]; // @[Shift.scala 66:70]
  assign _T_284 = _T_283[1]; // @[Shift.scala 12:21]
  assign _T_285 = _T_282[26:0]; // @[Shift.scala 64:52]
  assign _T_287 = {_T_285,2'h0}; // @[Cat.scala 29:58]
  assign _T_288 = _T_284 ? _T_287 : _T_282; // @[Shift.scala 64:27]
  assign _T_289 = _T_283[0:0]; // @[Shift.scala 66:70]
  assign _T_291 = _T_288[27:0]; // @[Shift.scala 64:52]
  assign _T_292 = {_T_291,1'h0}; // @[Cat.scala 29:58]
  assign _T_293 = _T_289 ? _T_292 : _T_288; // @[Shift.scala 64:27]
  assign _T_294 = _T_264 ? _T_293 : 29'h0; // @[Shift.scala 16:10]
  assign _T_295 = _T_294[28:28]; // @[convert.scala 23:34]
  assign decA_fraction = _T_294[27:0]; // @[convert.scala 24:34]
  assign _T_297 = _T_15 == 1'h0; // @[convert.scala 25:26]
  assign _T_299 = _T_15 ? _T_262 : _T_261; // @[convert.scala 25:42]
  assign _T_302 = ~ _T_295; // @[convert.scala 26:67]
  assign _T_303 = _T_13 ? _T_302 : _T_295; // @[convert.scala 26:51]
  assign _T_304 = {_T_297,_T_299,_T_303}; // @[Cat.scala 29:58]
  assign _T_306 = realA[30:0]; // @[convert.scala 29:56]
  assign _T_307 = _T_306 != 31'h0; // @[convert.scala 29:60]
  assign _T_308 = ~ _T_307; // @[convert.scala 29:41]
  assign decA_isNaR = _T_13 & _T_308; // @[convert.scala 29:39]
  assign _T_311 = _T_13 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_311 & _T_308; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_304); // @[convert.scala 32:24]
  assign _T_320 = io_B[31]; // @[convert.scala 18:24]
  assign _T_321 = io_B[30]; // @[convert.scala 18:40]
  assign _T_322 = _T_320 ^ _T_321; // @[convert.scala 18:36]
  assign _T_323 = io_B[30:1]; // @[convert.scala 19:24]
  assign _T_324 = io_B[29:0]; // @[convert.scala 19:43]
  assign _T_325 = _T_323 ^ _T_324; // @[convert.scala 19:39]
  assign _T_326 = _T_325[29:14]; // @[LZD.scala 43:32]
  assign _T_327 = _T_326[15:8]; // @[LZD.scala 43:32]
  assign _T_328 = _T_327[7:4]; // @[LZD.scala 43:32]
  assign _T_329 = _T_328[3:2]; // @[LZD.scala 43:32]
  assign _T_330 = _T_329 != 2'h0; // @[LZD.scala 39:14]
  assign _T_331 = _T_329[1]; // @[LZD.scala 39:21]
  assign _T_332 = _T_329[0]; // @[LZD.scala 39:30]
  assign _T_333 = ~ _T_332; // @[LZD.scala 39:27]
  assign _T_334 = _T_331 | _T_333; // @[LZD.scala 39:25]
  assign _T_335 = {_T_330,_T_334}; // @[Cat.scala 29:58]
  assign _T_336 = _T_328[1:0]; // @[LZD.scala 44:32]
  assign _T_337 = _T_336 != 2'h0; // @[LZD.scala 39:14]
  assign _T_338 = _T_336[1]; // @[LZD.scala 39:21]
  assign _T_339 = _T_336[0]; // @[LZD.scala 39:30]
  assign _T_340 = ~ _T_339; // @[LZD.scala 39:27]
  assign _T_341 = _T_338 | _T_340; // @[LZD.scala 39:25]
  assign _T_342 = {_T_337,_T_341}; // @[Cat.scala 29:58]
  assign _T_343 = _T_335[1]; // @[Shift.scala 12:21]
  assign _T_344 = _T_342[1]; // @[Shift.scala 12:21]
  assign _T_345 = _T_343 | _T_344; // @[LZD.scala 49:16]
  assign _T_346 = ~ _T_344; // @[LZD.scala 49:27]
  assign _T_347 = _T_343 | _T_346; // @[LZD.scala 49:25]
  assign _T_348 = _T_335[0:0]; // @[LZD.scala 49:47]
  assign _T_349 = _T_342[0:0]; // @[LZD.scala 49:59]
  assign _T_350 = _T_343 ? _T_348 : _T_349; // @[LZD.scala 49:35]
  assign _T_352 = {_T_345,_T_347,_T_350}; // @[Cat.scala 29:58]
  assign _T_353 = _T_327[3:0]; // @[LZD.scala 44:32]
  assign _T_354 = _T_353[3:2]; // @[LZD.scala 43:32]
  assign _T_355 = _T_354 != 2'h0; // @[LZD.scala 39:14]
  assign _T_356 = _T_354[1]; // @[LZD.scala 39:21]
  assign _T_357 = _T_354[0]; // @[LZD.scala 39:30]
  assign _T_358 = ~ _T_357; // @[LZD.scala 39:27]
  assign _T_359 = _T_356 | _T_358; // @[LZD.scala 39:25]
  assign _T_360 = {_T_355,_T_359}; // @[Cat.scala 29:58]
  assign _T_361 = _T_353[1:0]; // @[LZD.scala 44:32]
  assign _T_362 = _T_361 != 2'h0; // @[LZD.scala 39:14]
  assign _T_363 = _T_361[1]; // @[LZD.scala 39:21]
  assign _T_364 = _T_361[0]; // @[LZD.scala 39:30]
  assign _T_365 = ~ _T_364; // @[LZD.scala 39:27]
  assign _T_366 = _T_363 | _T_365; // @[LZD.scala 39:25]
  assign _T_367 = {_T_362,_T_366}; // @[Cat.scala 29:58]
  assign _T_368 = _T_360[1]; // @[Shift.scala 12:21]
  assign _T_369 = _T_367[1]; // @[Shift.scala 12:21]
  assign _T_370 = _T_368 | _T_369; // @[LZD.scala 49:16]
  assign _T_371 = ~ _T_369; // @[LZD.scala 49:27]
  assign _T_372 = _T_368 | _T_371; // @[LZD.scala 49:25]
  assign _T_373 = _T_360[0:0]; // @[LZD.scala 49:47]
  assign _T_374 = _T_367[0:0]; // @[LZD.scala 49:59]
  assign _T_375 = _T_368 ? _T_373 : _T_374; // @[LZD.scala 49:35]
  assign _T_377 = {_T_370,_T_372,_T_375}; // @[Cat.scala 29:58]
  assign _T_378 = _T_352[2]; // @[Shift.scala 12:21]
  assign _T_379 = _T_377[2]; // @[Shift.scala 12:21]
  assign _T_380 = _T_378 | _T_379; // @[LZD.scala 49:16]
  assign _T_381 = ~ _T_379; // @[LZD.scala 49:27]
  assign _T_382 = _T_378 | _T_381; // @[LZD.scala 49:25]
  assign _T_383 = _T_352[1:0]; // @[LZD.scala 49:47]
  assign _T_384 = _T_377[1:0]; // @[LZD.scala 49:59]
  assign _T_385 = _T_378 ? _T_383 : _T_384; // @[LZD.scala 49:35]
  assign _T_387 = {_T_380,_T_382,_T_385}; // @[Cat.scala 29:58]
  assign _T_388 = _T_326[7:0]; // @[LZD.scala 44:32]
  assign _T_389 = _T_388[7:4]; // @[LZD.scala 43:32]
  assign _T_390 = _T_389[3:2]; // @[LZD.scala 43:32]
  assign _T_391 = _T_390 != 2'h0; // @[LZD.scala 39:14]
  assign _T_392 = _T_390[1]; // @[LZD.scala 39:21]
  assign _T_393 = _T_390[0]; // @[LZD.scala 39:30]
  assign _T_394 = ~ _T_393; // @[LZD.scala 39:27]
  assign _T_395 = _T_392 | _T_394; // @[LZD.scala 39:25]
  assign _T_396 = {_T_391,_T_395}; // @[Cat.scala 29:58]
  assign _T_397 = _T_389[1:0]; // @[LZD.scala 44:32]
  assign _T_398 = _T_397 != 2'h0; // @[LZD.scala 39:14]
  assign _T_399 = _T_397[1]; // @[LZD.scala 39:21]
  assign _T_400 = _T_397[0]; // @[LZD.scala 39:30]
  assign _T_401 = ~ _T_400; // @[LZD.scala 39:27]
  assign _T_402 = _T_399 | _T_401; // @[LZD.scala 39:25]
  assign _T_403 = {_T_398,_T_402}; // @[Cat.scala 29:58]
  assign _T_404 = _T_396[1]; // @[Shift.scala 12:21]
  assign _T_405 = _T_403[1]; // @[Shift.scala 12:21]
  assign _T_406 = _T_404 | _T_405; // @[LZD.scala 49:16]
  assign _T_407 = ~ _T_405; // @[LZD.scala 49:27]
  assign _T_408 = _T_404 | _T_407; // @[LZD.scala 49:25]
  assign _T_409 = _T_396[0:0]; // @[LZD.scala 49:47]
  assign _T_410 = _T_403[0:0]; // @[LZD.scala 49:59]
  assign _T_411 = _T_404 ? _T_409 : _T_410; // @[LZD.scala 49:35]
  assign _T_413 = {_T_406,_T_408,_T_411}; // @[Cat.scala 29:58]
  assign _T_414 = _T_388[3:0]; // @[LZD.scala 44:32]
  assign _T_415 = _T_414[3:2]; // @[LZD.scala 43:32]
  assign _T_416 = _T_415 != 2'h0; // @[LZD.scala 39:14]
  assign _T_417 = _T_415[1]; // @[LZD.scala 39:21]
  assign _T_418 = _T_415[0]; // @[LZD.scala 39:30]
  assign _T_419 = ~ _T_418; // @[LZD.scala 39:27]
  assign _T_420 = _T_417 | _T_419; // @[LZD.scala 39:25]
  assign _T_421 = {_T_416,_T_420}; // @[Cat.scala 29:58]
  assign _T_422 = _T_414[1:0]; // @[LZD.scala 44:32]
  assign _T_423 = _T_422 != 2'h0; // @[LZD.scala 39:14]
  assign _T_424 = _T_422[1]; // @[LZD.scala 39:21]
  assign _T_425 = _T_422[0]; // @[LZD.scala 39:30]
  assign _T_426 = ~ _T_425; // @[LZD.scala 39:27]
  assign _T_427 = _T_424 | _T_426; // @[LZD.scala 39:25]
  assign _T_428 = {_T_423,_T_427}; // @[Cat.scala 29:58]
  assign _T_429 = _T_421[1]; // @[Shift.scala 12:21]
  assign _T_430 = _T_428[1]; // @[Shift.scala 12:21]
  assign _T_431 = _T_429 | _T_430; // @[LZD.scala 49:16]
  assign _T_432 = ~ _T_430; // @[LZD.scala 49:27]
  assign _T_433 = _T_429 | _T_432; // @[LZD.scala 49:25]
  assign _T_434 = _T_421[0:0]; // @[LZD.scala 49:47]
  assign _T_435 = _T_428[0:0]; // @[LZD.scala 49:59]
  assign _T_436 = _T_429 ? _T_434 : _T_435; // @[LZD.scala 49:35]
  assign _T_438 = {_T_431,_T_433,_T_436}; // @[Cat.scala 29:58]
  assign _T_439 = _T_413[2]; // @[Shift.scala 12:21]
  assign _T_440 = _T_438[2]; // @[Shift.scala 12:21]
  assign _T_441 = _T_439 | _T_440; // @[LZD.scala 49:16]
  assign _T_442 = ~ _T_440; // @[LZD.scala 49:27]
  assign _T_443 = _T_439 | _T_442; // @[LZD.scala 49:25]
  assign _T_444 = _T_413[1:0]; // @[LZD.scala 49:47]
  assign _T_445 = _T_438[1:0]; // @[LZD.scala 49:59]
  assign _T_446 = _T_439 ? _T_444 : _T_445; // @[LZD.scala 49:35]
  assign _T_448 = {_T_441,_T_443,_T_446}; // @[Cat.scala 29:58]
  assign _T_449 = _T_387[3]; // @[Shift.scala 12:21]
  assign _T_450 = _T_448[3]; // @[Shift.scala 12:21]
  assign _T_451 = _T_449 | _T_450; // @[LZD.scala 49:16]
  assign _T_452 = ~ _T_450; // @[LZD.scala 49:27]
  assign _T_453 = _T_449 | _T_452; // @[LZD.scala 49:25]
  assign _T_454 = _T_387[2:0]; // @[LZD.scala 49:47]
  assign _T_455 = _T_448[2:0]; // @[LZD.scala 49:59]
  assign _T_456 = _T_449 ? _T_454 : _T_455; // @[LZD.scala 49:35]
  assign _T_458 = {_T_451,_T_453,_T_456}; // @[Cat.scala 29:58]
  assign _T_459 = _T_325[13:0]; // @[LZD.scala 44:32]
  assign _T_460 = _T_459[13:6]; // @[LZD.scala 43:32]
  assign _T_461 = _T_460[7:4]; // @[LZD.scala 43:32]
  assign _T_462 = _T_461[3:2]; // @[LZD.scala 43:32]
  assign _T_463 = _T_462 != 2'h0; // @[LZD.scala 39:14]
  assign _T_464 = _T_462[1]; // @[LZD.scala 39:21]
  assign _T_465 = _T_462[0]; // @[LZD.scala 39:30]
  assign _T_466 = ~ _T_465; // @[LZD.scala 39:27]
  assign _T_467 = _T_464 | _T_466; // @[LZD.scala 39:25]
  assign _T_468 = {_T_463,_T_467}; // @[Cat.scala 29:58]
  assign _T_469 = _T_461[1:0]; // @[LZD.scala 44:32]
  assign _T_470 = _T_469 != 2'h0; // @[LZD.scala 39:14]
  assign _T_471 = _T_469[1]; // @[LZD.scala 39:21]
  assign _T_472 = _T_469[0]; // @[LZD.scala 39:30]
  assign _T_473 = ~ _T_472; // @[LZD.scala 39:27]
  assign _T_474 = _T_471 | _T_473; // @[LZD.scala 39:25]
  assign _T_475 = {_T_470,_T_474}; // @[Cat.scala 29:58]
  assign _T_476 = _T_468[1]; // @[Shift.scala 12:21]
  assign _T_477 = _T_475[1]; // @[Shift.scala 12:21]
  assign _T_478 = _T_476 | _T_477; // @[LZD.scala 49:16]
  assign _T_479 = ~ _T_477; // @[LZD.scala 49:27]
  assign _T_480 = _T_476 | _T_479; // @[LZD.scala 49:25]
  assign _T_481 = _T_468[0:0]; // @[LZD.scala 49:47]
  assign _T_482 = _T_475[0:0]; // @[LZD.scala 49:59]
  assign _T_483 = _T_476 ? _T_481 : _T_482; // @[LZD.scala 49:35]
  assign _T_485 = {_T_478,_T_480,_T_483}; // @[Cat.scala 29:58]
  assign _T_486 = _T_460[3:0]; // @[LZD.scala 44:32]
  assign _T_487 = _T_486[3:2]; // @[LZD.scala 43:32]
  assign _T_488 = _T_487 != 2'h0; // @[LZD.scala 39:14]
  assign _T_489 = _T_487[1]; // @[LZD.scala 39:21]
  assign _T_490 = _T_487[0]; // @[LZD.scala 39:30]
  assign _T_491 = ~ _T_490; // @[LZD.scala 39:27]
  assign _T_492 = _T_489 | _T_491; // @[LZD.scala 39:25]
  assign _T_493 = {_T_488,_T_492}; // @[Cat.scala 29:58]
  assign _T_494 = _T_486[1:0]; // @[LZD.scala 44:32]
  assign _T_495 = _T_494 != 2'h0; // @[LZD.scala 39:14]
  assign _T_496 = _T_494[1]; // @[LZD.scala 39:21]
  assign _T_497 = _T_494[0]; // @[LZD.scala 39:30]
  assign _T_498 = ~ _T_497; // @[LZD.scala 39:27]
  assign _T_499 = _T_496 | _T_498; // @[LZD.scala 39:25]
  assign _T_500 = {_T_495,_T_499}; // @[Cat.scala 29:58]
  assign _T_501 = _T_493[1]; // @[Shift.scala 12:21]
  assign _T_502 = _T_500[1]; // @[Shift.scala 12:21]
  assign _T_503 = _T_501 | _T_502; // @[LZD.scala 49:16]
  assign _T_504 = ~ _T_502; // @[LZD.scala 49:27]
  assign _T_505 = _T_501 | _T_504; // @[LZD.scala 49:25]
  assign _T_506 = _T_493[0:0]; // @[LZD.scala 49:47]
  assign _T_507 = _T_500[0:0]; // @[LZD.scala 49:59]
  assign _T_508 = _T_501 ? _T_506 : _T_507; // @[LZD.scala 49:35]
  assign _T_510 = {_T_503,_T_505,_T_508}; // @[Cat.scala 29:58]
  assign _T_511 = _T_485[2]; // @[Shift.scala 12:21]
  assign _T_512 = _T_510[2]; // @[Shift.scala 12:21]
  assign _T_513 = _T_511 | _T_512; // @[LZD.scala 49:16]
  assign _T_514 = ~ _T_512; // @[LZD.scala 49:27]
  assign _T_515 = _T_511 | _T_514; // @[LZD.scala 49:25]
  assign _T_516 = _T_485[1:0]; // @[LZD.scala 49:47]
  assign _T_517 = _T_510[1:0]; // @[LZD.scala 49:59]
  assign _T_518 = _T_511 ? _T_516 : _T_517; // @[LZD.scala 49:35]
  assign _T_520 = {_T_513,_T_515,_T_518}; // @[Cat.scala 29:58]
  assign _T_521 = _T_459[5:0]; // @[LZD.scala 44:32]
  assign _T_522 = _T_521[5:2]; // @[LZD.scala 43:32]
  assign _T_523 = _T_522[3:2]; // @[LZD.scala 43:32]
  assign _T_524 = _T_523 != 2'h0; // @[LZD.scala 39:14]
  assign _T_525 = _T_523[1]; // @[LZD.scala 39:21]
  assign _T_526 = _T_523[0]; // @[LZD.scala 39:30]
  assign _T_527 = ~ _T_526; // @[LZD.scala 39:27]
  assign _T_528 = _T_525 | _T_527; // @[LZD.scala 39:25]
  assign _T_529 = {_T_524,_T_528}; // @[Cat.scala 29:58]
  assign _T_530 = _T_522[1:0]; // @[LZD.scala 44:32]
  assign _T_531 = _T_530 != 2'h0; // @[LZD.scala 39:14]
  assign _T_532 = _T_530[1]; // @[LZD.scala 39:21]
  assign _T_533 = _T_530[0]; // @[LZD.scala 39:30]
  assign _T_534 = ~ _T_533; // @[LZD.scala 39:27]
  assign _T_535 = _T_532 | _T_534; // @[LZD.scala 39:25]
  assign _T_536 = {_T_531,_T_535}; // @[Cat.scala 29:58]
  assign _T_537 = _T_529[1]; // @[Shift.scala 12:21]
  assign _T_538 = _T_536[1]; // @[Shift.scala 12:21]
  assign _T_539 = _T_537 | _T_538; // @[LZD.scala 49:16]
  assign _T_540 = ~ _T_538; // @[LZD.scala 49:27]
  assign _T_541 = _T_537 | _T_540; // @[LZD.scala 49:25]
  assign _T_542 = _T_529[0:0]; // @[LZD.scala 49:47]
  assign _T_543 = _T_536[0:0]; // @[LZD.scala 49:59]
  assign _T_544 = _T_537 ? _T_542 : _T_543; // @[LZD.scala 49:35]
  assign _T_546 = {_T_539,_T_541,_T_544}; // @[Cat.scala 29:58]
  assign _T_547 = _T_521[1:0]; // @[LZD.scala 44:32]
  assign _T_548 = _T_547 != 2'h0; // @[LZD.scala 39:14]
  assign _T_549 = _T_547[1]; // @[LZD.scala 39:21]
  assign _T_550 = _T_547[0]; // @[LZD.scala 39:30]
  assign _T_551 = ~ _T_550; // @[LZD.scala 39:27]
  assign _T_552 = _T_549 | _T_551; // @[LZD.scala 39:25]
  assign _T_553 = {_T_548,_T_552}; // @[Cat.scala 29:58]
  assign _T_554 = _T_546[2]; // @[Shift.scala 12:21]
  assign _T_556 = _T_546[1:0]; // @[LZD.scala 55:32]
  assign _T_557 = _T_554 ? _T_556 : _T_553; // @[LZD.scala 55:20]
  assign _T_558 = {_T_554,_T_557}; // @[Cat.scala 29:58]
  assign _T_559 = _T_520[3]; // @[Shift.scala 12:21]
  assign _T_561 = _T_520[2:0]; // @[LZD.scala 55:32]
  assign _T_562 = _T_559 ? _T_561 : _T_558; // @[LZD.scala 55:20]
  assign _T_563 = {_T_559,_T_562}; // @[Cat.scala 29:58]
  assign _T_564 = _T_458[4]; // @[Shift.scala 12:21]
  assign _T_566 = _T_458[3:0]; // @[LZD.scala 55:32]
  assign _T_567 = _T_564 ? _T_566 : _T_563; // @[LZD.scala 55:20]
  assign _T_568 = {_T_564,_T_567}; // @[Cat.scala 29:58]
  assign _T_569 = ~ _T_568; // @[convert.scala 21:22]
  assign _T_570 = io_B[28:0]; // @[convert.scala 22:36]
  assign _T_571 = _T_569 < 5'h1d; // @[Shift.scala 16:24]
  assign _T_573 = _T_569[4]; // @[Shift.scala 12:21]
  assign _T_574 = _T_570[12:0]; // @[Shift.scala 64:52]
  assign _T_576 = {_T_574,16'h0}; // @[Cat.scala 29:58]
  assign _T_577 = _T_573 ? _T_576 : _T_570; // @[Shift.scala 64:27]
  assign _T_578 = _T_569[3:0]; // @[Shift.scala 66:70]
  assign _T_579 = _T_578[3]; // @[Shift.scala 12:21]
  assign _T_580 = _T_577[20:0]; // @[Shift.scala 64:52]
  assign _T_582 = {_T_580,8'h0}; // @[Cat.scala 29:58]
  assign _T_583 = _T_579 ? _T_582 : _T_577; // @[Shift.scala 64:27]
  assign _T_584 = _T_578[2:0]; // @[Shift.scala 66:70]
  assign _T_585 = _T_584[2]; // @[Shift.scala 12:21]
  assign _T_586 = _T_583[24:0]; // @[Shift.scala 64:52]
  assign _T_588 = {_T_586,4'h0}; // @[Cat.scala 29:58]
  assign _T_589 = _T_585 ? _T_588 : _T_583; // @[Shift.scala 64:27]
  assign _T_590 = _T_584[1:0]; // @[Shift.scala 66:70]
  assign _T_591 = _T_590[1]; // @[Shift.scala 12:21]
  assign _T_592 = _T_589[26:0]; // @[Shift.scala 64:52]
  assign _T_594 = {_T_592,2'h0}; // @[Cat.scala 29:58]
  assign _T_595 = _T_591 ? _T_594 : _T_589; // @[Shift.scala 64:27]
  assign _T_596 = _T_590[0:0]; // @[Shift.scala 66:70]
  assign _T_598 = _T_595[27:0]; // @[Shift.scala 64:52]
  assign _T_599 = {_T_598,1'h0}; // @[Cat.scala 29:58]
  assign _T_600 = _T_596 ? _T_599 : _T_595; // @[Shift.scala 64:27]
  assign _T_601 = _T_571 ? _T_600 : 29'h0; // @[Shift.scala 16:10]
  assign _T_602 = _T_601[28:28]; // @[convert.scala 23:34]
  assign decB_fraction = _T_601[27:0]; // @[convert.scala 24:34]
  assign _T_604 = _T_322 == 1'h0; // @[convert.scala 25:26]
  assign _T_606 = _T_322 ? _T_569 : _T_568; // @[convert.scala 25:42]
  assign _T_609 = ~ _T_602; // @[convert.scala 26:67]
  assign _T_610 = _T_320 ? _T_609 : _T_602; // @[convert.scala 26:51]
  assign _T_611 = {_T_604,_T_606,_T_610}; // @[Cat.scala 29:58]
  assign _T_613 = io_B[30:0]; // @[convert.scala 29:56]
  assign _T_614 = _T_613 != 31'h0; // @[convert.scala 29:60]
  assign _T_615 = ~ _T_614; // @[convert.scala 29:41]
  assign decB_isNaR = _T_320 & _T_615; // @[convert.scala 29:39]
  assign _T_618 = _T_320 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_618 & _T_615; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_611); // @[convert.scala 32:24]
  assign _T_627 = realC[31]; // @[convert.scala 18:24]
  assign _T_628 = realC[30]; // @[convert.scala 18:40]
  assign _T_629 = _T_627 ^ _T_628; // @[convert.scala 18:36]
  assign _T_630 = realC[30:1]; // @[convert.scala 19:24]
  assign _T_631 = realC[29:0]; // @[convert.scala 19:43]
  assign _T_632 = _T_630 ^ _T_631; // @[convert.scala 19:39]
  assign _T_633 = _T_632[29:14]; // @[LZD.scala 43:32]
  assign _T_634 = _T_633[15:8]; // @[LZD.scala 43:32]
  assign _T_635 = _T_634[7:4]; // @[LZD.scala 43:32]
  assign _T_636 = _T_635[3:2]; // @[LZD.scala 43:32]
  assign _T_637 = _T_636 != 2'h0; // @[LZD.scala 39:14]
  assign _T_638 = _T_636[1]; // @[LZD.scala 39:21]
  assign _T_639 = _T_636[0]; // @[LZD.scala 39:30]
  assign _T_640 = ~ _T_639; // @[LZD.scala 39:27]
  assign _T_641 = _T_638 | _T_640; // @[LZD.scala 39:25]
  assign _T_642 = {_T_637,_T_641}; // @[Cat.scala 29:58]
  assign _T_643 = _T_635[1:0]; // @[LZD.scala 44:32]
  assign _T_644 = _T_643 != 2'h0; // @[LZD.scala 39:14]
  assign _T_645 = _T_643[1]; // @[LZD.scala 39:21]
  assign _T_646 = _T_643[0]; // @[LZD.scala 39:30]
  assign _T_647 = ~ _T_646; // @[LZD.scala 39:27]
  assign _T_648 = _T_645 | _T_647; // @[LZD.scala 39:25]
  assign _T_649 = {_T_644,_T_648}; // @[Cat.scala 29:58]
  assign _T_650 = _T_642[1]; // @[Shift.scala 12:21]
  assign _T_651 = _T_649[1]; // @[Shift.scala 12:21]
  assign _T_652 = _T_650 | _T_651; // @[LZD.scala 49:16]
  assign _T_653 = ~ _T_651; // @[LZD.scala 49:27]
  assign _T_654 = _T_650 | _T_653; // @[LZD.scala 49:25]
  assign _T_655 = _T_642[0:0]; // @[LZD.scala 49:47]
  assign _T_656 = _T_649[0:0]; // @[LZD.scala 49:59]
  assign _T_657 = _T_650 ? _T_655 : _T_656; // @[LZD.scala 49:35]
  assign _T_659 = {_T_652,_T_654,_T_657}; // @[Cat.scala 29:58]
  assign _T_660 = _T_634[3:0]; // @[LZD.scala 44:32]
  assign _T_661 = _T_660[3:2]; // @[LZD.scala 43:32]
  assign _T_662 = _T_661 != 2'h0; // @[LZD.scala 39:14]
  assign _T_663 = _T_661[1]; // @[LZD.scala 39:21]
  assign _T_664 = _T_661[0]; // @[LZD.scala 39:30]
  assign _T_665 = ~ _T_664; // @[LZD.scala 39:27]
  assign _T_666 = _T_663 | _T_665; // @[LZD.scala 39:25]
  assign _T_667 = {_T_662,_T_666}; // @[Cat.scala 29:58]
  assign _T_668 = _T_660[1:0]; // @[LZD.scala 44:32]
  assign _T_669 = _T_668 != 2'h0; // @[LZD.scala 39:14]
  assign _T_670 = _T_668[1]; // @[LZD.scala 39:21]
  assign _T_671 = _T_668[0]; // @[LZD.scala 39:30]
  assign _T_672 = ~ _T_671; // @[LZD.scala 39:27]
  assign _T_673 = _T_670 | _T_672; // @[LZD.scala 39:25]
  assign _T_674 = {_T_669,_T_673}; // @[Cat.scala 29:58]
  assign _T_675 = _T_667[1]; // @[Shift.scala 12:21]
  assign _T_676 = _T_674[1]; // @[Shift.scala 12:21]
  assign _T_677 = _T_675 | _T_676; // @[LZD.scala 49:16]
  assign _T_678 = ~ _T_676; // @[LZD.scala 49:27]
  assign _T_679 = _T_675 | _T_678; // @[LZD.scala 49:25]
  assign _T_680 = _T_667[0:0]; // @[LZD.scala 49:47]
  assign _T_681 = _T_674[0:0]; // @[LZD.scala 49:59]
  assign _T_682 = _T_675 ? _T_680 : _T_681; // @[LZD.scala 49:35]
  assign _T_684 = {_T_677,_T_679,_T_682}; // @[Cat.scala 29:58]
  assign _T_685 = _T_659[2]; // @[Shift.scala 12:21]
  assign _T_686 = _T_684[2]; // @[Shift.scala 12:21]
  assign _T_687 = _T_685 | _T_686; // @[LZD.scala 49:16]
  assign _T_688 = ~ _T_686; // @[LZD.scala 49:27]
  assign _T_689 = _T_685 | _T_688; // @[LZD.scala 49:25]
  assign _T_690 = _T_659[1:0]; // @[LZD.scala 49:47]
  assign _T_691 = _T_684[1:0]; // @[LZD.scala 49:59]
  assign _T_692 = _T_685 ? _T_690 : _T_691; // @[LZD.scala 49:35]
  assign _T_694 = {_T_687,_T_689,_T_692}; // @[Cat.scala 29:58]
  assign _T_695 = _T_633[7:0]; // @[LZD.scala 44:32]
  assign _T_696 = _T_695[7:4]; // @[LZD.scala 43:32]
  assign _T_697 = _T_696[3:2]; // @[LZD.scala 43:32]
  assign _T_698 = _T_697 != 2'h0; // @[LZD.scala 39:14]
  assign _T_699 = _T_697[1]; // @[LZD.scala 39:21]
  assign _T_700 = _T_697[0]; // @[LZD.scala 39:30]
  assign _T_701 = ~ _T_700; // @[LZD.scala 39:27]
  assign _T_702 = _T_699 | _T_701; // @[LZD.scala 39:25]
  assign _T_703 = {_T_698,_T_702}; // @[Cat.scala 29:58]
  assign _T_704 = _T_696[1:0]; // @[LZD.scala 44:32]
  assign _T_705 = _T_704 != 2'h0; // @[LZD.scala 39:14]
  assign _T_706 = _T_704[1]; // @[LZD.scala 39:21]
  assign _T_707 = _T_704[0]; // @[LZD.scala 39:30]
  assign _T_708 = ~ _T_707; // @[LZD.scala 39:27]
  assign _T_709 = _T_706 | _T_708; // @[LZD.scala 39:25]
  assign _T_710 = {_T_705,_T_709}; // @[Cat.scala 29:58]
  assign _T_711 = _T_703[1]; // @[Shift.scala 12:21]
  assign _T_712 = _T_710[1]; // @[Shift.scala 12:21]
  assign _T_713 = _T_711 | _T_712; // @[LZD.scala 49:16]
  assign _T_714 = ~ _T_712; // @[LZD.scala 49:27]
  assign _T_715 = _T_711 | _T_714; // @[LZD.scala 49:25]
  assign _T_716 = _T_703[0:0]; // @[LZD.scala 49:47]
  assign _T_717 = _T_710[0:0]; // @[LZD.scala 49:59]
  assign _T_718 = _T_711 ? _T_716 : _T_717; // @[LZD.scala 49:35]
  assign _T_720 = {_T_713,_T_715,_T_718}; // @[Cat.scala 29:58]
  assign _T_721 = _T_695[3:0]; // @[LZD.scala 44:32]
  assign _T_722 = _T_721[3:2]; // @[LZD.scala 43:32]
  assign _T_723 = _T_722 != 2'h0; // @[LZD.scala 39:14]
  assign _T_724 = _T_722[1]; // @[LZD.scala 39:21]
  assign _T_725 = _T_722[0]; // @[LZD.scala 39:30]
  assign _T_726 = ~ _T_725; // @[LZD.scala 39:27]
  assign _T_727 = _T_724 | _T_726; // @[LZD.scala 39:25]
  assign _T_728 = {_T_723,_T_727}; // @[Cat.scala 29:58]
  assign _T_729 = _T_721[1:0]; // @[LZD.scala 44:32]
  assign _T_730 = _T_729 != 2'h0; // @[LZD.scala 39:14]
  assign _T_731 = _T_729[1]; // @[LZD.scala 39:21]
  assign _T_732 = _T_729[0]; // @[LZD.scala 39:30]
  assign _T_733 = ~ _T_732; // @[LZD.scala 39:27]
  assign _T_734 = _T_731 | _T_733; // @[LZD.scala 39:25]
  assign _T_735 = {_T_730,_T_734}; // @[Cat.scala 29:58]
  assign _T_736 = _T_728[1]; // @[Shift.scala 12:21]
  assign _T_737 = _T_735[1]; // @[Shift.scala 12:21]
  assign _T_738 = _T_736 | _T_737; // @[LZD.scala 49:16]
  assign _T_739 = ~ _T_737; // @[LZD.scala 49:27]
  assign _T_740 = _T_736 | _T_739; // @[LZD.scala 49:25]
  assign _T_741 = _T_728[0:0]; // @[LZD.scala 49:47]
  assign _T_742 = _T_735[0:0]; // @[LZD.scala 49:59]
  assign _T_743 = _T_736 ? _T_741 : _T_742; // @[LZD.scala 49:35]
  assign _T_745 = {_T_738,_T_740,_T_743}; // @[Cat.scala 29:58]
  assign _T_746 = _T_720[2]; // @[Shift.scala 12:21]
  assign _T_747 = _T_745[2]; // @[Shift.scala 12:21]
  assign _T_748 = _T_746 | _T_747; // @[LZD.scala 49:16]
  assign _T_749 = ~ _T_747; // @[LZD.scala 49:27]
  assign _T_750 = _T_746 | _T_749; // @[LZD.scala 49:25]
  assign _T_751 = _T_720[1:0]; // @[LZD.scala 49:47]
  assign _T_752 = _T_745[1:0]; // @[LZD.scala 49:59]
  assign _T_753 = _T_746 ? _T_751 : _T_752; // @[LZD.scala 49:35]
  assign _T_755 = {_T_748,_T_750,_T_753}; // @[Cat.scala 29:58]
  assign _T_756 = _T_694[3]; // @[Shift.scala 12:21]
  assign _T_757 = _T_755[3]; // @[Shift.scala 12:21]
  assign _T_758 = _T_756 | _T_757; // @[LZD.scala 49:16]
  assign _T_759 = ~ _T_757; // @[LZD.scala 49:27]
  assign _T_760 = _T_756 | _T_759; // @[LZD.scala 49:25]
  assign _T_761 = _T_694[2:0]; // @[LZD.scala 49:47]
  assign _T_762 = _T_755[2:0]; // @[LZD.scala 49:59]
  assign _T_763 = _T_756 ? _T_761 : _T_762; // @[LZD.scala 49:35]
  assign _T_765 = {_T_758,_T_760,_T_763}; // @[Cat.scala 29:58]
  assign _T_766 = _T_632[13:0]; // @[LZD.scala 44:32]
  assign _T_767 = _T_766[13:6]; // @[LZD.scala 43:32]
  assign _T_768 = _T_767[7:4]; // @[LZD.scala 43:32]
  assign _T_769 = _T_768[3:2]; // @[LZD.scala 43:32]
  assign _T_770 = _T_769 != 2'h0; // @[LZD.scala 39:14]
  assign _T_771 = _T_769[1]; // @[LZD.scala 39:21]
  assign _T_772 = _T_769[0]; // @[LZD.scala 39:30]
  assign _T_773 = ~ _T_772; // @[LZD.scala 39:27]
  assign _T_774 = _T_771 | _T_773; // @[LZD.scala 39:25]
  assign _T_775 = {_T_770,_T_774}; // @[Cat.scala 29:58]
  assign _T_776 = _T_768[1:0]; // @[LZD.scala 44:32]
  assign _T_777 = _T_776 != 2'h0; // @[LZD.scala 39:14]
  assign _T_778 = _T_776[1]; // @[LZD.scala 39:21]
  assign _T_779 = _T_776[0]; // @[LZD.scala 39:30]
  assign _T_780 = ~ _T_779; // @[LZD.scala 39:27]
  assign _T_781 = _T_778 | _T_780; // @[LZD.scala 39:25]
  assign _T_782 = {_T_777,_T_781}; // @[Cat.scala 29:58]
  assign _T_783 = _T_775[1]; // @[Shift.scala 12:21]
  assign _T_784 = _T_782[1]; // @[Shift.scala 12:21]
  assign _T_785 = _T_783 | _T_784; // @[LZD.scala 49:16]
  assign _T_786 = ~ _T_784; // @[LZD.scala 49:27]
  assign _T_787 = _T_783 | _T_786; // @[LZD.scala 49:25]
  assign _T_788 = _T_775[0:0]; // @[LZD.scala 49:47]
  assign _T_789 = _T_782[0:0]; // @[LZD.scala 49:59]
  assign _T_790 = _T_783 ? _T_788 : _T_789; // @[LZD.scala 49:35]
  assign _T_792 = {_T_785,_T_787,_T_790}; // @[Cat.scala 29:58]
  assign _T_793 = _T_767[3:0]; // @[LZD.scala 44:32]
  assign _T_794 = _T_793[3:2]; // @[LZD.scala 43:32]
  assign _T_795 = _T_794 != 2'h0; // @[LZD.scala 39:14]
  assign _T_796 = _T_794[1]; // @[LZD.scala 39:21]
  assign _T_797 = _T_794[0]; // @[LZD.scala 39:30]
  assign _T_798 = ~ _T_797; // @[LZD.scala 39:27]
  assign _T_799 = _T_796 | _T_798; // @[LZD.scala 39:25]
  assign _T_800 = {_T_795,_T_799}; // @[Cat.scala 29:58]
  assign _T_801 = _T_793[1:0]; // @[LZD.scala 44:32]
  assign _T_802 = _T_801 != 2'h0; // @[LZD.scala 39:14]
  assign _T_803 = _T_801[1]; // @[LZD.scala 39:21]
  assign _T_804 = _T_801[0]; // @[LZD.scala 39:30]
  assign _T_805 = ~ _T_804; // @[LZD.scala 39:27]
  assign _T_806 = _T_803 | _T_805; // @[LZD.scala 39:25]
  assign _T_807 = {_T_802,_T_806}; // @[Cat.scala 29:58]
  assign _T_808 = _T_800[1]; // @[Shift.scala 12:21]
  assign _T_809 = _T_807[1]; // @[Shift.scala 12:21]
  assign _T_810 = _T_808 | _T_809; // @[LZD.scala 49:16]
  assign _T_811 = ~ _T_809; // @[LZD.scala 49:27]
  assign _T_812 = _T_808 | _T_811; // @[LZD.scala 49:25]
  assign _T_813 = _T_800[0:0]; // @[LZD.scala 49:47]
  assign _T_814 = _T_807[0:0]; // @[LZD.scala 49:59]
  assign _T_815 = _T_808 ? _T_813 : _T_814; // @[LZD.scala 49:35]
  assign _T_817 = {_T_810,_T_812,_T_815}; // @[Cat.scala 29:58]
  assign _T_818 = _T_792[2]; // @[Shift.scala 12:21]
  assign _T_819 = _T_817[2]; // @[Shift.scala 12:21]
  assign _T_820 = _T_818 | _T_819; // @[LZD.scala 49:16]
  assign _T_821 = ~ _T_819; // @[LZD.scala 49:27]
  assign _T_822 = _T_818 | _T_821; // @[LZD.scala 49:25]
  assign _T_823 = _T_792[1:0]; // @[LZD.scala 49:47]
  assign _T_824 = _T_817[1:0]; // @[LZD.scala 49:59]
  assign _T_825 = _T_818 ? _T_823 : _T_824; // @[LZD.scala 49:35]
  assign _T_827 = {_T_820,_T_822,_T_825}; // @[Cat.scala 29:58]
  assign _T_828 = _T_766[5:0]; // @[LZD.scala 44:32]
  assign _T_829 = _T_828[5:2]; // @[LZD.scala 43:32]
  assign _T_830 = _T_829[3:2]; // @[LZD.scala 43:32]
  assign _T_831 = _T_830 != 2'h0; // @[LZD.scala 39:14]
  assign _T_832 = _T_830[1]; // @[LZD.scala 39:21]
  assign _T_833 = _T_830[0]; // @[LZD.scala 39:30]
  assign _T_834 = ~ _T_833; // @[LZD.scala 39:27]
  assign _T_835 = _T_832 | _T_834; // @[LZD.scala 39:25]
  assign _T_836 = {_T_831,_T_835}; // @[Cat.scala 29:58]
  assign _T_837 = _T_829[1:0]; // @[LZD.scala 44:32]
  assign _T_838 = _T_837 != 2'h0; // @[LZD.scala 39:14]
  assign _T_839 = _T_837[1]; // @[LZD.scala 39:21]
  assign _T_840 = _T_837[0]; // @[LZD.scala 39:30]
  assign _T_841 = ~ _T_840; // @[LZD.scala 39:27]
  assign _T_842 = _T_839 | _T_841; // @[LZD.scala 39:25]
  assign _T_843 = {_T_838,_T_842}; // @[Cat.scala 29:58]
  assign _T_844 = _T_836[1]; // @[Shift.scala 12:21]
  assign _T_845 = _T_843[1]; // @[Shift.scala 12:21]
  assign _T_846 = _T_844 | _T_845; // @[LZD.scala 49:16]
  assign _T_847 = ~ _T_845; // @[LZD.scala 49:27]
  assign _T_848 = _T_844 | _T_847; // @[LZD.scala 49:25]
  assign _T_849 = _T_836[0:0]; // @[LZD.scala 49:47]
  assign _T_850 = _T_843[0:0]; // @[LZD.scala 49:59]
  assign _T_851 = _T_844 ? _T_849 : _T_850; // @[LZD.scala 49:35]
  assign _T_853 = {_T_846,_T_848,_T_851}; // @[Cat.scala 29:58]
  assign _T_854 = _T_828[1:0]; // @[LZD.scala 44:32]
  assign _T_855 = _T_854 != 2'h0; // @[LZD.scala 39:14]
  assign _T_856 = _T_854[1]; // @[LZD.scala 39:21]
  assign _T_857 = _T_854[0]; // @[LZD.scala 39:30]
  assign _T_858 = ~ _T_857; // @[LZD.scala 39:27]
  assign _T_859 = _T_856 | _T_858; // @[LZD.scala 39:25]
  assign _T_860 = {_T_855,_T_859}; // @[Cat.scala 29:58]
  assign _T_861 = _T_853[2]; // @[Shift.scala 12:21]
  assign _T_863 = _T_853[1:0]; // @[LZD.scala 55:32]
  assign _T_864 = _T_861 ? _T_863 : _T_860; // @[LZD.scala 55:20]
  assign _T_865 = {_T_861,_T_864}; // @[Cat.scala 29:58]
  assign _T_866 = _T_827[3]; // @[Shift.scala 12:21]
  assign _T_868 = _T_827[2:0]; // @[LZD.scala 55:32]
  assign _T_869 = _T_866 ? _T_868 : _T_865; // @[LZD.scala 55:20]
  assign _T_870 = {_T_866,_T_869}; // @[Cat.scala 29:58]
  assign _T_871 = _T_765[4]; // @[Shift.scala 12:21]
  assign _T_873 = _T_765[3:0]; // @[LZD.scala 55:32]
  assign _T_874 = _T_871 ? _T_873 : _T_870; // @[LZD.scala 55:20]
  assign _T_875 = {_T_871,_T_874}; // @[Cat.scala 29:58]
  assign _T_876 = ~ _T_875; // @[convert.scala 21:22]
  assign _T_877 = realC[28:0]; // @[convert.scala 22:36]
  assign _T_878 = _T_876 < 5'h1d; // @[Shift.scala 16:24]
  assign _T_880 = _T_876[4]; // @[Shift.scala 12:21]
  assign _T_881 = _T_877[12:0]; // @[Shift.scala 64:52]
  assign _T_883 = {_T_881,16'h0}; // @[Cat.scala 29:58]
  assign _T_884 = _T_880 ? _T_883 : _T_877; // @[Shift.scala 64:27]
  assign _T_885 = _T_876[3:0]; // @[Shift.scala 66:70]
  assign _T_886 = _T_885[3]; // @[Shift.scala 12:21]
  assign _T_887 = _T_884[20:0]; // @[Shift.scala 64:52]
  assign _T_889 = {_T_887,8'h0}; // @[Cat.scala 29:58]
  assign _T_890 = _T_886 ? _T_889 : _T_884; // @[Shift.scala 64:27]
  assign _T_891 = _T_885[2:0]; // @[Shift.scala 66:70]
  assign _T_892 = _T_891[2]; // @[Shift.scala 12:21]
  assign _T_893 = _T_890[24:0]; // @[Shift.scala 64:52]
  assign _T_895 = {_T_893,4'h0}; // @[Cat.scala 29:58]
  assign _T_896 = _T_892 ? _T_895 : _T_890; // @[Shift.scala 64:27]
  assign _T_897 = _T_891[1:0]; // @[Shift.scala 66:70]
  assign _T_898 = _T_897[1]; // @[Shift.scala 12:21]
  assign _T_899 = _T_896[26:0]; // @[Shift.scala 64:52]
  assign _T_901 = {_T_899,2'h0}; // @[Cat.scala 29:58]
  assign _T_902 = _T_898 ? _T_901 : _T_896; // @[Shift.scala 64:27]
  assign _T_903 = _T_897[0:0]; // @[Shift.scala 66:70]
  assign _T_905 = _T_902[27:0]; // @[Shift.scala 64:52]
  assign _T_906 = {_T_905,1'h0}; // @[Cat.scala 29:58]
  assign _T_907 = _T_903 ? _T_906 : _T_902; // @[Shift.scala 64:27]
  assign _T_908 = _T_878 ? _T_907 : 29'h0; // @[Shift.scala 16:10]
  assign _T_909 = _T_908[28:28]; // @[convert.scala 23:34]
  assign decC_fraction = _T_908[27:0]; // @[convert.scala 24:34]
  assign _T_911 = _T_629 == 1'h0; // @[convert.scala 25:26]
  assign _T_913 = _T_629 ? _T_876 : _T_875; // @[convert.scala 25:42]
  assign _T_916 = ~ _T_909; // @[convert.scala 26:67]
  assign _T_917 = _T_627 ? _T_916 : _T_909; // @[convert.scala 26:51]
  assign _T_918 = {_T_911,_T_913,_T_917}; // @[Cat.scala 29:58]
  assign _T_920 = realC[30:0]; // @[convert.scala 29:56]
  assign _T_921 = _T_920 != 31'h0; // @[convert.scala 29:60]
  assign _T_922 = ~ _T_921; // @[convert.scala 29:41]
  assign decC_isNaR = _T_627 & _T_922; // @[convert.scala 29:39]
  assign _T_925 = _T_627 == 1'h0; // @[convert.scala 30:19]
  assign decC_isZero = _T_925 & _T_922; // @[convert.scala 30:41]
  assign decC_scale = $signed(_T_918); // @[convert.scala 32:24]
  assign _T_933 = decA_isNaR | decB_isNaR; // @[PositFMA.scala 58:30]
  assign outIsNaR = _T_933 | decC_isNaR; // @[PositFMA.scala 58:44]
  assign _T_934 = ~ _T_13; // @[PositFMA.scala 59:34]
  assign _T_935 = ~ decA_isZero; // @[PositFMA.scala 59:47]
  assign _T_936 = _T_934 & _T_935; // @[PositFMA.scala 59:45]
  assign _T_938 = {_T_13,_T_936,decA_fraction}; // @[Cat.scala 29:58]
  assign sigA = $signed(_T_938); // @[PositFMA.scala 59:76]
  assign _T_939 = ~ _T_320; // @[PositFMA.scala 60:34]
  assign _T_940 = ~ decB_isZero; // @[PositFMA.scala 60:47]
  assign _T_941 = _T_939 & _T_940; // @[PositFMA.scala 60:45]
  assign _T_943 = {_T_320,_T_941,decB_fraction}; // @[Cat.scala 29:58]
  assign sigB = $signed(_T_943); // @[PositFMA.scala 60:76]
  assign _T_944 = $signed(sigA) * $signed(sigB); // @[PositFMA.scala 61:25]
  assign sigP = $unsigned(_T_944); // @[PositFMA.scala 61:33]
  assign head2 = sigP[59:58]; // @[PositFMA.scala 62:28]
  assign _T_945 = head2[1]; // @[PositFMA.scala 63:31]
  assign _T_946 = ~ _T_945; // @[PositFMA.scala 63:25]
  assign _T_947 = head2[0]; // @[PositFMA.scala 63:42]
  assign addTwo = _T_946 & _T_947; // @[PositFMA.scala 63:35]
  assign _T_948 = sigP[59]; // @[PositFMA.scala 65:23]
  assign _T_949 = sigP[57]; // @[PositFMA.scala 65:49]
  assign addOne = _T_948 ^ _T_949; // @[PositFMA.scala 65:43]
  assign _T_950 = {addTwo,addOne}; // @[Cat.scala 29:58]
  assign expBias = {1'b0,$signed(_T_950)}; // @[PositFMA.scala 66:39]
  assign mulSign = sigP[59:59]; // @[PositFMA.scala 67:28]
  assign _T_951 = $signed(decA_scale) + $signed(decB_scale); // @[PositFMA.scala 69:30]
  assign _GEN_12 = {{5{expBias[2]}},expBias}; // @[PositFMA.scala 69:44]
  assign _T_953 = $signed(_T_951) + $signed(_GEN_12); // @[PositFMA.scala 69:44]
  assign mulScale = $signed(_T_953); // @[PositFMA.scala 69:44]
  assign _T_954 = sigP[57:0]; // @[PositFMA.scala 72:29]
  assign _T_955 = sigP[56:0]; // @[PositFMA.scala 73:29]
  assign _T_956 = {_T_955, 1'h0}; // @[PositFMA.scala 73:48]
  assign mulSigTmp = addOne ? _T_954 : _T_956; // @[PositFMA.scala 70:22]
  assign _T_958 = mulSigTmp[57:57]; // @[PositFMA.scala 77:39]
  assign _T_959 = _T_958 | addTwo; // @[PositFMA.scala 77:43]
  assign _T_960 = mulSigTmp[56:0]; // @[PositFMA.scala 78:39]
  assign mulSig = {mulSign,_T_959,_T_960}; // @[Cat.scala 29:58]
  assign _T_986 = ~ addSign_phase2; // @[PositFMA.scala 107:29]
  assign _T_987 = ~ addZero_phase2; // @[PositFMA.scala 107:47]
  assign _T_988 = _T_986 & _T_987; // @[PositFMA.scala 107:45]
  assign extAddSig = {addSign_phase2,_T_988,addFrac_phase2,29'h0}; // @[Cat.scala 29:58]
  assign _GEN_13 = {{1{addScale_phase2[6]}},addScale_phase2}; // @[PositFMA.scala 111:39]
  assign mulGreater = $signed(mulScale_phase2) > $signed(_GEN_13); // @[PositFMA.scala 111:39]
  assign greaterScale = mulGreater ? $signed(mulScale_phase2) : $signed({{1{addScale_phase2[6]}},addScale_phase2}); // @[PositFMA.scala 112:26]
  assign smallerScale = mulGreater ? $signed({{1{addScale_phase2[6]}},addScale_phase2}) : $signed(mulScale_phase2); // @[PositFMA.scala 113:26]
  assign _T_992 = $signed(greaterScale) - $signed(smallerScale); // @[PositFMA.scala 114:36]
  assign scaleDiff = $signed(_T_992); // @[PositFMA.scala 114:36]
  assign greaterSig = mulGreater ? mulSig_phase2 : extAddSig; // @[PositFMA.scala 115:26]
  assign smallerSigTmp = mulGreater ? extAddSig : mulSig_phase2; // @[PositFMA.scala 116:26]
  assign _T_993 = $unsigned(scaleDiff); // @[PositFMA.scala 117:69]
  assign _T_994 = _T_993 < 8'h3b; // @[Shift.scala 39:24]
  assign _T_995 = _T_993[5:0]; // @[Shift.scala 40:44]
  assign _T_996 = smallerSigTmp[58:32]; // @[Shift.scala 90:30]
  assign _T_997 = smallerSigTmp[31:0]; // @[Shift.scala 90:48]
  assign _T_998 = _T_997 != 32'h0; // @[Shift.scala 90:57]
  assign _GEN_14 = {{26'd0}, _T_998}; // @[Shift.scala 90:39]
  assign _T_999 = _T_996 | _GEN_14; // @[Shift.scala 90:39]
  assign _T_1000 = _T_995[5]; // @[Shift.scala 12:21]
  assign _T_1001 = smallerSigTmp[58]; // @[Shift.scala 12:21]
  assign _T_1003 = _T_1001 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 71:12]
  assign _T_1004 = {_T_1003,_T_999}; // @[Cat.scala 29:58]
  assign _T_1005 = _T_1000 ? _T_1004 : smallerSigTmp; // @[Shift.scala 91:22]
  assign _T_1006 = _T_995[4:0]; // @[Shift.scala 92:77]
  assign _T_1007 = _T_1005[58:16]; // @[Shift.scala 90:30]
  assign _T_1008 = _T_1005[15:0]; // @[Shift.scala 90:48]
  assign _T_1009 = _T_1008 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_15 = {{42'd0}, _T_1009}; // @[Shift.scala 90:39]
  assign _T_1010 = _T_1007 | _GEN_15; // @[Shift.scala 90:39]
  assign _T_1011 = _T_1006[4]; // @[Shift.scala 12:21]
  assign _T_1012 = _T_1005[58]; // @[Shift.scala 12:21]
  assign _T_1014 = _T_1012 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_1015 = {_T_1014,_T_1010}; // @[Cat.scala 29:58]
  assign _T_1016 = _T_1011 ? _T_1015 : _T_1005; // @[Shift.scala 91:22]
  assign _T_1017 = _T_1006[3:0]; // @[Shift.scala 92:77]
  assign _T_1018 = _T_1016[58:8]; // @[Shift.scala 90:30]
  assign _T_1019 = _T_1016[7:0]; // @[Shift.scala 90:48]
  assign _T_1020 = _T_1019 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_16 = {{50'd0}, _T_1020}; // @[Shift.scala 90:39]
  assign _T_1021 = _T_1018 | _GEN_16; // @[Shift.scala 90:39]
  assign _T_1022 = _T_1017[3]; // @[Shift.scala 12:21]
  assign _T_1023 = _T_1016[58]; // @[Shift.scala 12:21]
  assign _T_1025 = _T_1023 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_1026 = {_T_1025,_T_1021}; // @[Cat.scala 29:58]
  assign _T_1027 = _T_1022 ? _T_1026 : _T_1016; // @[Shift.scala 91:22]
  assign _T_1028 = _T_1017[2:0]; // @[Shift.scala 92:77]
  assign _T_1029 = _T_1027[58:4]; // @[Shift.scala 90:30]
  assign _T_1030 = _T_1027[3:0]; // @[Shift.scala 90:48]
  assign _T_1031 = _T_1030 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_17 = {{54'd0}, _T_1031}; // @[Shift.scala 90:39]
  assign _T_1032 = _T_1029 | _GEN_17; // @[Shift.scala 90:39]
  assign _T_1033 = _T_1028[2]; // @[Shift.scala 12:21]
  assign _T_1034 = _T_1027[58]; // @[Shift.scala 12:21]
  assign _T_1036 = _T_1034 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_1037 = {_T_1036,_T_1032}; // @[Cat.scala 29:58]
  assign _T_1038 = _T_1033 ? _T_1037 : _T_1027; // @[Shift.scala 91:22]
  assign _T_1039 = _T_1028[1:0]; // @[Shift.scala 92:77]
  assign _T_1040 = _T_1038[58:2]; // @[Shift.scala 90:30]
  assign _T_1041 = _T_1038[1:0]; // @[Shift.scala 90:48]
  assign _T_1042 = _T_1041 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_18 = {{56'd0}, _T_1042}; // @[Shift.scala 90:39]
  assign _T_1043 = _T_1040 | _GEN_18; // @[Shift.scala 90:39]
  assign _T_1044 = _T_1039[1]; // @[Shift.scala 12:21]
  assign _T_1045 = _T_1038[58]; // @[Shift.scala 12:21]
  assign _T_1047 = _T_1045 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_1048 = {_T_1047,_T_1043}; // @[Cat.scala 29:58]
  assign _T_1049 = _T_1044 ? _T_1048 : _T_1038; // @[Shift.scala 91:22]
  assign _T_1050 = _T_1039[0:0]; // @[Shift.scala 92:77]
  assign _T_1051 = _T_1049[58:1]; // @[Shift.scala 90:30]
  assign _T_1052 = _T_1049[0:0]; // @[Shift.scala 90:48]
  assign _GEN_19 = {{57'd0}, _T_1052}; // @[Shift.scala 90:39]
  assign _T_1054 = _T_1051 | _GEN_19; // @[Shift.scala 90:39]
  assign _T_1056 = _T_1049[58]; // @[Shift.scala 12:21]
  assign _T_1057 = {_T_1056,_T_1054}; // @[Cat.scala 29:58]
  assign _T_1058 = _T_1050 ? _T_1057 : _T_1049; // @[Shift.scala 91:22]
  assign _T_1061 = _T_1001 ? 59'h7ffffffffffffff : 59'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_994 ? _T_1058 : _T_1061; // @[Shift.scala 39:10]
  assign rawSumSig = greaterSig + smallerSig; // @[PositFMA.scala 118:34]
  assign _T_1062 = mulSig_phase2[58:58]; // @[PositFMA.scala 119:42]
  assign _T_1063 = _T_1062 ^ addSign_phase2; // @[PositFMA.scala 119:46]
  assign _T_1064 = rawSumSig[59:59]; // @[PositFMA.scala 119:79]
  assign sumSign = _T_1063 ^ _T_1064; // @[PositFMA.scala 119:63]
  assign _T_1066 = greaterSig + smallerSig; // @[PositFMA.scala 120:50]
  assign signSumSig = {sumSign,_T_1066}; // @[Cat.scala 29:58]
  assign _T_1067 = signSumSig[59:1]; // @[PositFMA.scala 124:33]
  assign _T_1068 = signSumSig[58:0]; // @[PositFMA.scala 124:68]
  assign sumXor = _T_1067 ^ _T_1068; // @[PositFMA.scala 124:51]
  assign _T_1069 = sumXor[58:27]; // @[LZD.scala 43:32]
  assign _T_1070 = _T_1069[31:16]; // @[LZD.scala 43:32]
  assign _T_1071 = _T_1070[15:8]; // @[LZD.scala 43:32]
  assign _T_1072 = _T_1071[7:4]; // @[LZD.scala 43:32]
  assign _T_1073 = _T_1072[3:2]; // @[LZD.scala 43:32]
  assign _T_1074 = _T_1073 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1075 = _T_1073[1]; // @[LZD.scala 39:21]
  assign _T_1076 = _T_1073[0]; // @[LZD.scala 39:30]
  assign _T_1077 = ~ _T_1076; // @[LZD.scala 39:27]
  assign _T_1078 = _T_1075 | _T_1077; // @[LZD.scala 39:25]
  assign _T_1079 = {_T_1074,_T_1078}; // @[Cat.scala 29:58]
  assign _T_1080 = _T_1072[1:0]; // @[LZD.scala 44:32]
  assign _T_1081 = _T_1080 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1082 = _T_1080[1]; // @[LZD.scala 39:21]
  assign _T_1083 = _T_1080[0]; // @[LZD.scala 39:30]
  assign _T_1084 = ~ _T_1083; // @[LZD.scala 39:27]
  assign _T_1085 = _T_1082 | _T_1084; // @[LZD.scala 39:25]
  assign _T_1086 = {_T_1081,_T_1085}; // @[Cat.scala 29:58]
  assign _T_1087 = _T_1079[1]; // @[Shift.scala 12:21]
  assign _T_1088 = _T_1086[1]; // @[Shift.scala 12:21]
  assign _T_1089 = _T_1087 | _T_1088; // @[LZD.scala 49:16]
  assign _T_1090 = ~ _T_1088; // @[LZD.scala 49:27]
  assign _T_1091 = _T_1087 | _T_1090; // @[LZD.scala 49:25]
  assign _T_1092 = _T_1079[0:0]; // @[LZD.scala 49:47]
  assign _T_1093 = _T_1086[0:0]; // @[LZD.scala 49:59]
  assign _T_1094 = _T_1087 ? _T_1092 : _T_1093; // @[LZD.scala 49:35]
  assign _T_1096 = {_T_1089,_T_1091,_T_1094}; // @[Cat.scala 29:58]
  assign _T_1097 = _T_1071[3:0]; // @[LZD.scala 44:32]
  assign _T_1098 = _T_1097[3:2]; // @[LZD.scala 43:32]
  assign _T_1099 = _T_1098 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1100 = _T_1098[1]; // @[LZD.scala 39:21]
  assign _T_1101 = _T_1098[0]; // @[LZD.scala 39:30]
  assign _T_1102 = ~ _T_1101; // @[LZD.scala 39:27]
  assign _T_1103 = _T_1100 | _T_1102; // @[LZD.scala 39:25]
  assign _T_1104 = {_T_1099,_T_1103}; // @[Cat.scala 29:58]
  assign _T_1105 = _T_1097[1:0]; // @[LZD.scala 44:32]
  assign _T_1106 = _T_1105 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1107 = _T_1105[1]; // @[LZD.scala 39:21]
  assign _T_1108 = _T_1105[0]; // @[LZD.scala 39:30]
  assign _T_1109 = ~ _T_1108; // @[LZD.scala 39:27]
  assign _T_1110 = _T_1107 | _T_1109; // @[LZD.scala 39:25]
  assign _T_1111 = {_T_1106,_T_1110}; // @[Cat.scala 29:58]
  assign _T_1112 = _T_1104[1]; // @[Shift.scala 12:21]
  assign _T_1113 = _T_1111[1]; // @[Shift.scala 12:21]
  assign _T_1114 = _T_1112 | _T_1113; // @[LZD.scala 49:16]
  assign _T_1115 = ~ _T_1113; // @[LZD.scala 49:27]
  assign _T_1116 = _T_1112 | _T_1115; // @[LZD.scala 49:25]
  assign _T_1117 = _T_1104[0:0]; // @[LZD.scala 49:47]
  assign _T_1118 = _T_1111[0:0]; // @[LZD.scala 49:59]
  assign _T_1119 = _T_1112 ? _T_1117 : _T_1118; // @[LZD.scala 49:35]
  assign _T_1121 = {_T_1114,_T_1116,_T_1119}; // @[Cat.scala 29:58]
  assign _T_1122 = _T_1096[2]; // @[Shift.scala 12:21]
  assign _T_1123 = _T_1121[2]; // @[Shift.scala 12:21]
  assign _T_1124 = _T_1122 | _T_1123; // @[LZD.scala 49:16]
  assign _T_1125 = ~ _T_1123; // @[LZD.scala 49:27]
  assign _T_1126 = _T_1122 | _T_1125; // @[LZD.scala 49:25]
  assign _T_1127 = _T_1096[1:0]; // @[LZD.scala 49:47]
  assign _T_1128 = _T_1121[1:0]; // @[LZD.scala 49:59]
  assign _T_1129 = _T_1122 ? _T_1127 : _T_1128; // @[LZD.scala 49:35]
  assign _T_1131 = {_T_1124,_T_1126,_T_1129}; // @[Cat.scala 29:58]
  assign _T_1132 = _T_1070[7:0]; // @[LZD.scala 44:32]
  assign _T_1133 = _T_1132[7:4]; // @[LZD.scala 43:32]
  assign _T_1134 = _T_1133[3:2]; // @[LZD.scala 43:32]
  assign _T_1135 = _T_1134 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1136 = _T_1134[1]; // @[LZD.scala 39:21]
  assign _T_1137 = _T_1134[0]; // @[LZD.scala 39:30]
  assign _T_1138 = ~ _T_1137; // @[LZD.scala 39:27]
  assign _T_1139 = _T_1136 | _T_1138; // @[LZD.scala 39:25]
  assign _T_1140 = {_T_1135,_T_1139}; // @[Cat.scala 29:58]
  assign _T_1141 = _T_1133[1:0]; // @[LZD.scala 44:32]
  assign _T_1142 = _T_1141 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1143 = _T_1141[1]; // @[LZD.scala 39:21]
  assign _T_1144 = _T_1141[0]; // @[LZD.scala 39:30]
  assign _T_1145 = ~ _T_1144; // @[LZD.scala 39:27]
  assign _T_1146 = _T_1143 | _T_1145; // @[LZD.scala 39:25]
  assign _T_1147 = {_T_1142,_T_1146}; // @[Cat.scala 29:58]
  assign _T_1148 = _T_1140[1]; // @[Shift.scala 12:21]
  assign _T_1149 = _T_1147[1]; // @[Shift.scala 12:21]
  assign _T_1150 = _T_1148 | _T_1149; // @[LZD.scala 49:16]
  assign _T_1151 = ~ _T_1149; // @[LZD.scala 49:27]
  assign _T_1152 = _T_1148 | _T_1151; // @[LZD.scala 49:25]
  assign _T_1153 = _T_1140[0:0]; // @[LZD.scala 49:47]
  assign _T_1154 = _T_1147[0:0]; // @[LZD.scala 49:59]
  assign _T_1155 = _T_1148 ? _T_1153 : _T_1154; // @[LZD.scala 49:35]
  assign _T_1157 = {_T_1150,_T_1152,_T_1155}; // @[Cat.scala 29:58]
  assign _T_1158 = _T_1132[3:0]; // @[LZD.scala 44:32]
  assign _T_1159 = _T_1158[3:2]; // @[LZD.scala 43:32]
  assign _T_1160 = _T_1159 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1161 = _T_1159[1]; // @[LZD.scala 39:21]
  assign _T_1162 = _T_1159[0]; // @[LZD.scala 39:30]
  assign _T_1163 = ~ _T_1162; // @[LZD.scala 39:27]
  assign _T_1164 = _T_1161 | _T_1163; // @[LZD.scala 39:25]
  assign _T_1165 = {_T_1160,_T_1164}; // @[Cat.scala 29:58]
  assign _T_1166 = _T_1158[1:0]; // @[LZD.scala 44:32]
  assign _T_1167 = _T_1166 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1168 = _T_1166[1]; // @[LZD.scala 39:21]
  assign _T_1169 = _T_1166[0]; // @[LZD.scala 39:30]
  assign _T_1170 = ~ _T_1169; // @[LZD.scala 39:27]
  assign _T_1171 = _T_1168 | _T_1170; // @[LZD.scala 39:25]
  assign _T_1172 = {_T_1167,_T_1171}; // @[Cat.scala 29:58]
  assign _T_1173 = _T_1165[1]; // @[Shift.scala 12:21]
  assign _T_1174 = _T_1172[1]; // @[Shift.scala 12:21]
  assign _T_1175 = _T_1173 | _T_1174; // @[LZD.scala 49:16]
  assign _T_1176 = ~ _T_1174; // @[LZD.scala 49:27]
  assign _T_1177 = _T_1173 | _T_1176; // @[LZD.scala 49:25]
  assign _T_1178 = _T_1165[0:0]; // @[LZD.scala 49:47]
  assign _T_1179 = _T_1172[0:0]; // @[LZD.scala 49:59]
  assign _T_1180 = _T_1173 ? _T_1178 : _T_1179; // @[LZD.scala 49:35]
  assign _T_1182 = {_T_1175,_T_1177,_T_1180}; // @[Cat.scala 29:58]
  assign _T_1183 = _T_1157[2]; // @[Shift.scala 12:21]
  assign _T_1184 = _T_1182[2]; // @[Shift.scala 12:21]
  assign _T_1185 = _T_1183 | _T_1184; // @[LZD.scala 49:16]
  assign _T_1186 = ~ _T_1184; // @[LZD.scala 49:27]
  assign _T_1187 = _T_1183 | _T_1186; // @[LZD.scala 49:25]
  assign _T_1188 = _T_1157[1:0]; // @[LZD.scala 49:47]
  assign _T_1189 = _T_1182[1:0]; // @[LZD.scala 49:59]
  assign _T_1190 = _T_1183 ? _T_1188 : _T_1189; // @[LZD.scala 49:35]
  assign _T_1192 = {_T_1185,_T_1187,_T_1190}; // @[Cat.scala 29:58]
  assign _T_1193 = _T_1131[3]; // @[Shift.scala 12:21]
  assign _T_1194 = _T_1192[3]; // @[Shift.scala 12:21]
  assign _T_1195 = _T_1193 | _T_1194; // @[LZD.scala 49:16]
  assign _T_1196 = ~ _T_1194; // @[LZD.scala 49:27]
  assign _T_1197 = _T_1193 | _T_1196; // @[LZD.scala 49:25]
  assign _T_1198 = _T_1131[2:0]; // @[LZD.scala 49:47]
  assign _T_1199 = _T_1192[2:0]; // @[LZD.scala 49:59]
  assign _T_1200 = _T_1193 ? _T_1198 : _T_1199; // @[LZD.scala 49:35]
  assign _T_1202 = {_T_1195,_T_1197,_T_1200}; // @[Cat.scala 29:58]
  assign _T_1203 = _T_1069[15:0]; // @[LZD.scala 44:32]
  assign _T_1204 = _T_1203[15:8]; // @[LZD.scala 43:32]
  assign _T_1205 = _T_1204[7:4]; // @[LZD.scala 43:32]
  assign _T_1206 = _T_1205[3:2]; // @[LZD.scala 43:32]
  assign _T_1207 = _T_1206 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1208 = _T_1206[1]; // @[LZD.scala 39:21]
  assign _T_1209 = _T_1206[0]; // @[LZD.scala 39:30]
  assign _T_1210 = ~ _T_1209; // @[LZD.scala 39:27]
  assign _T_1211 = _T_1208 | _T_1210; // @[LZD.scala 39:25]
  assign _T_1212 = {_T_1207,_T_1211}; // @[Cat.scala 29:58]
  assign _T_1213 = _T_1205[1:0]; // @[LZD.scala 44:32]
  assign _T_1214 = _T_1213 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1215 = _T_1213[1]; // @[LZD.scala 39:21]
  assign _T_1216 = _T_1213[0]; // @[LZD.scala 39:30]
  assign _T_1217 = ~ _T_1216; // @[LZD.scala 39:27]
  assign _T_1218 = _T_1215 | _T_1217; // @[LZD.scala 39:25]
  assign _T_1219 = {_T_1214,_T_1218}; // @[Cat.scala 29:58]
  assign _T_1220 = _T_1212[1]; // @[Shift.scala 12:21]
  assign _T_1221 = _T_1219[1]; // @[Shift.scala 12:21]
  assign _T_1222 = _T_1220 | _T_1221; // @[LZD.scala 49:16]
  assign _T_1223 = ~ _T_1221; // @[LZD.scala 49:27]
  assign _T_1224 = _T_1220 | _T_1223; // @[LZD.scala 49:25]
  assign _T_1225 = _T_1212[0:0]; // @[LZD.scala 49:47]
  assign _T_1226 = _T_1219[0:0]; // @[LZD.scala 49:59]
  assign _T_1227 = _T_1220 ? _T_1225 : _T_1226; // @[LZD.scala 49:35]
  assign _T_1229 = {_T_1222,_T_1224,_T_1227}; // @[Cat.scala 29:58]
  assign _T_1230 = _T_1204[3:0]; // @[LZD.scala 44:32]
  assign _T_1231 = _T_1230[3:2]; // @[LZD.scala 43:32]
  assign _T_1232 = _T_1231 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1233 = _T_1231[1]; // @[LZD.scala 39:21]
  assign _T_1234 = _T_1231[0]; // @[LZD.scala 39:30]
  assign _T_1235 = ~ _T_1234; // @[LZD.scala 39:27]
  assign _T_1236 = _T_1233 | _T_1235; // @[LZD.scala 39:25]
  assign _T_1237 = {_T_1232,_T_1236}; // @[Cat.scala 29:58]
  assign _T_1238 = _T_1230[1:0]; // @[LZD.scala 44:32]
  assign _T_1239 = _T_1238 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1240 = _T_1238[1]; // @[LZD.scala 39:21]
  assign _T_1241 = _T_1238[0]; // @[LZD.scala 39:30]
  assign _T_1242 = ~ _T_1241; // @[LZD.scala 39:27]
  assign _T_1243 = _T_1240 | _T_1242; // @[LZD.scala 39:25]
  assign _T_1244 = {_T_1239,_T_1243}; // @[Cat.scala 29:58]
  assign _T_1245 = _T_1237[1]; // @[Shift.scala 12:21]
  assign _T_1246 = _T_1244[1]; // @[Shift.scala 12:21]
  assign _T_1247 = _T_1245 | _T_1246; // @[LZD.scala 49:16]
  assign _T_1248 = ~ _T_1246; // @[LZD.scala 49:27]
  assign _T_1249 = _T_1245 | _T_1248; // @[LZD.scala 49:25]
  assign _T_1250 = _T_1237[0:0]; // @[LZD.scala 49:47]
  assign _T_1251 = _T_1244[0:0]; // @[LZD.scala 49:59]
  assign _T_1252 = _T_1245 ? _T_1250 : _T_1251; // @[LZD.scala 49:35]
  assign _T_1254 = {_T_1247,_T_1249,_T_1252}; // @[Cat.scala 29:58]
  assign _T_1255 = _T_1229[2]; // @[Shift.scala 12:21]
  assign _T_1256 = _T_1254[2]; // @[Shift.scala 12:21]
  assign _T_1257 = _T_1255 | _T_1256; // @[LZD.scala 49:16]
  assign _T_1258 = ~ _T_1256; // @[LZD.scala 49:27]
  assign _T_1259 = _T_1255 | _T_1258; // @[LZD.scala 49:25]
  assign _T_1260 = _T_1229[1:0]; // @[LZD.scala 49:47]
  assign _T_1261 = _T_1254[1:0]; // @[LZD.scala 49:59]
  assign _T_1262 = _T_1255 ? _T_1260 : _T_1261; // @[LZD.scala 49:35]
  assign _T_1264 = {_T_1257,_T_1259,_T_1262}; // @[Cat.scala 29:58]
  assign _T_1265 = _T_1203[7:0]; // @[LZD.scala 44:32]
  assign _T_1266 = _T_1265[7:4]; // @[LZD.scala 43:32]
  assign _T_1267 = _T_1266[3:2]; // @[LZD.scala 43:32]
  assign _T_1268 = _T_1267 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1269 = _T_1267[1]; // @[LZD.scala 39:21]
  assign _T_1270 = _T_1267[0]; // @[LZD.scala 39:30]
  assign _T_1271 = ~ _T_1270; // @[LZD.scala 39:27]
  assign _T_1272 = _T_1269 | _T_1271; // @[LZD.scala 39:25]
  assign _T_1273 = {_T_1268,_T_1272}; // @[Cat.scala 29:58]
  assign _T_1274 = _T_1266[1:0]; // @[LZD.scala 44:32]
  assign _T_1275 = _T_1274 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1276 = _T_1274[1]; // @[LZD.scala 39:21]
  assign _T_1277 = _T_1274[0]; // @[LZD.scala 39:30]
  assign _T_1278 = ~ _T_1277; // @[LZD.scala 39:27]
  assign _T_1279 = _T_1276 | _T_1278; // @[LZD.scala 39:25]
  assign _T_1280 = {_T_1275,_T_1279}; // @[Cat.scala 29:58]
  assign _T_1281 = _T_1273[1]; // @[Shift.scala 12:21]
  assign _T_1282 = _T_1280[1]; // @[Shift.scala 12:21]
  assign _T_1283 = _T_1281 | _T_1282; // @[LZD.scala 49:16]
  assign _T_1284 = ~ _T_1282; // @[LZD.scala 49:27]
  assign _T_1285 = _T_1281 | _T_1284; // @[LZD.scala 49:25]
  assign _T_1286 = _T_1273[0:0]; // @[LZD.scala 49:47]
  assign _T_1287 = _T_1280[0:0]; // @[LZD.scala 49:59]
  assign _T_1288 = _T_1281 ? _T_1286 : _T_1287; // @[LZD.scala 49:35]
  assign _T_1290 = {_T_1283,_T_1285,_T_1288}; // @[Cat.scala 29:58]
  assign _T_1291 = _T_1265[3:0]; // @[LZD.scala 44:32]
  assign _T_1292 = _T_1291[3:2]; // @[LZD.scala 43:32]
  assign _T_1293 = _T_1292 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1294 = _T_1292[1]; // @[LZD.scala 39:21]
  assign _T_1295 = _T_1292[0]; // @[LZD.scala 39:30]
  assign _T_1296 = ~ _T_1295; // @[LZD.scala 39:27]
  assign _T_1297 = _T_1294 | _T_1296; // @[LZD.scala 39:25]
  assign _T_1298 = {_T_1293,_T_1297}; // @[Cat.scala 29:58]
  assign _T_1299 = _T_1291[1:0]; // @[LZD.scala 44:32]
  assign _T_1300 = _T_1299 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1301 = _T_1299[1]; // @[LZD.scala 39:21]
  assign _T_1302 = _T_1299[0]; // @[LZD.scala 39:30]
  assign _T_1303 = ~ _T_1302; // @[LZD.scala 39:27]
  assign _T_1304 = _T_1301 | _T_1303; // @[LZD.scala 39:25]
  assign _T_1305 = {_T_1300,_T_1304}; // @[Cat.scala 29:58]
  assign _T_1306 = _T_1298[1]; // @[Shift.scala 12:21]
  assign _T_1307 = _T_1305[1]; // @[Shift.scala 12:21]
  assign _T_1308 = _T_1306 | _T_1307; // @[LZD.scala 49:16]
  assign _T_1309 = ~ _T_1307; // @[LZD.scala 49:27]
  assign _T_1310 = _T_1306 | _T_1309; // @[LZD.scala 49:25]
  assign _T_1311 = _T_1298[0:0]; // @[LZD.scala 49:47]
  assign _T_1312 = _T_1305[0:0]; // @[LZD.scala 49:59]
  assign _T_1313 = _T_1306 ? _T_1311 : _T_1312; // @[LZD.scala 49:35]
  assign _T_1315 = {_T_1308,_T_1310,_T_1313}; // @[Cat.scala 29:58]
  assign _T_1316 = _T_1290[2]; // @[Shift.scala 12:21]
  assign _T_1317 = _T_1315[2]; // @[Shift.scala 12:21]
  assign _T_1318 = _T_1316 | _T_1317; // @[LZD.scala 49:16]
  assign _T_1319 = ~ _T_1317; // @[LZD.scala 49:27]
  assign _T_1320 = _T_1316 | _T_1319; // @[LZD.scala 49:25]
  assign _T_1321 = _T_1290[1:0]; // @[LZD.scala 49:47]
  assign _T_1322 = _T_1315[1:0]; // @[LZD.scala 49:59]
  assign _T_1323 = _T_1316 ? _T_1321 : _T_1322; // @[LZD.scala 49:35]
  assign _T_1325 = {_T_1318,_T_1320,_T_1323}; // @[Cat.scala 29:58]
  assign _T_1326 = _T_1264[3]; // @[Shift.scala 12:21]
  assign _T_1327 = _T_1325[3]; // @[Shift.scala 12:21]
  assign _T_1328 = _T_1326 | _T_1327; // @[LZD.scala 49:16]
  assign _T_1329 = ~ _T_1327; // @[LZD.scala 49:27]
  assign _T_1330 = _T_1326 | _T_1329; // @[LZD.scala 49:25]
  assign _T_1331 = _T_1264[2:0]; // @[LZD.scala 49:47]
  assign _T_1332 = _T_1325[2:0]; // @[LZD.scala 49:59]
  assign _T_1333 = _T_1326 ? _T_1331 : _T_1332; // @[LZD.scala 49:35]
  assign _T_1335 = {_T_1328,_T_1330,_T_1333}; // @[Cat.scala 29:58]
  assign _T_1336 = _T_1202[4]; // @[Shift.scala 12:21]
  assign _T_1337 = _T_1335[4]; // @[Shift.scala 12:21]
  assign _T_1338 = _T_1336 | _T_1337; // @[LZD.scala 49:16]
  assign _T_1339 = ~ _T_1337; // @[LZD.scala 49:27]
  assign _T_1340 = _T_1336 | _T_1339; // @[LZD.scala 49:25]
  assign _T_1341 = _T_1202[3:0]; // @[LZD.scala 49:47]
  assign _T_1342 = _T_1335[3:0]; // @[LZD.scala 49:59]
  assign _T_1343 = _T_1336 ? _T_1341 : _T_1342; // @[LZD.scala 49:35]
  assign _T_1345 = {_T_1338,_T_1340,_T_1343}; // @[Cat.scala 29:58]
  assign _T_1346 = sumXor[26:0]; // @[LZD.scala 44:32]
  assign _T_1347 = _T_1346[26:11]; // @[LZD.scala 43:32]
  assign _T_1348 = _T_1347[15:8]; // @[LZD.scala 43:32]
  assign _T_1349 = _T_1348[7:4]; // @[LZD.scala 43:32]
  assign _T_1350 = _T_1349[3:2]; // @[LZD.scala 43:32]
  assign _T_1351 = _T_1350 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1352 = _T_1350[1]; // @[LZD.scala 39:21]
  assign _T_1353 = _T_1350[0]; // @[LZD.scala 39:30]
  assign _T_1354 = ~ _T_1353; // @[LZD.scala 39:27]
  assign _T_1355 = _T_1352 | _T_1354; // @[LZD.scala 39:25]
  assign _T_1356 = {_T_1351,_T_1355}; // @[Cat.scala 29:58]
  assign _T_1357 = _T_1349[1:0]; // @[LZD.scala 44:32]
  assign _T_1358 = _T_1357 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1359 = _T_1357[1]; // @[LZD.scala 39:21]
  assign _T_1360 = _T_1357[0]; // @[LZD.scala 39:30]
  assign _T_1361 = ~ _T_1360; // @[LZD.scala 39:27]
  assign _T_1362 = _T_1359 | _T_1361; // @[LZD.scala 39:25]
  assign _T_1363 = {_T_1358,_T_1362}; // @[Cat.scala 29:58]
  assign _T_1364 = _T_1356[1]; // @[Shift.scala 12:21]
  assign _T_1365 = _T_1363[1]; // @[Shift.scala 12:21]
  assign _T_1366 = _T_1364 | _T_1365; // @[LZD.scala 49:16]
  assign _T_1367 = ~ _T_1365; // @[LZD.scala 49:27]
  assign _T_1368 = _T_1364 | _T_1367; // @[LZD.scala 49:25]
  assign _T_1369 = _T_1356[0:0]; // @[LZD.scala 49:47]
  assign _T_1370 = _T_1363[0:0]; // @[LZD.scala 49:59]
  assign _T_1371 = _T_1364 ? _T_1369 : _T_1370; // @[LZD.scala 49:35]
  assign _T_1373 = {_T_1366,_T_1368,_T_1371}; // @[Cat.scala 29:58]
  assign _T_1374 = _T_1348[3:0]; // @[LZD.scala 44:32]
  assign _T_1375 = _T_1374[3:2]; // @[LZD.scala 43:32]
  assign _T_1376 = _T_1375 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1377 = _T_1375[1]; // @[LZD.scala 39:21]
  assign _T_1378 = _T_1375[0]; // @[LZD.scala 39:30]
  assign _T_1379 = ~ _T_1378; // @[LZD.scala 39:27]
  assign _T_1380 = _T_1377 | _T_1379; // @[LZD.scala 39:25]
  assign _T_1381 = {_T_1376,_T_1380}; // @[Cat.scala 29:58]
  assign _T_1382 = _T_1374[1:0]; // @[LZD.scala 44:32]
  assign _T_1383 = _T_1382 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1384 = _T_1382[1]; // @[LZD.scala 39:21]
  assign _T_1385 = _T_1382[0]; // @[LZD.scala 39:30]
  assign _T_1386 = ~ _T_1385; // @[LZD.scala 39:27]
  assign _T_1387 = _T_1384 | _T_1386; // @[LZD.scala 39:25]
  assign _T_1388 = {_T_1383,_T_1387}; // @[Cat.scala 29:58]
  assign _T_1389 = _T_1381[1]; // @[Shift.scala 12:21]
  assign _T_1390 = _T_1388[1]; // @[Shift.scala 12:21]
  assign _T_1391 = _T_1389 | _T_1390; // @[LZD.scala 49:16]
  assign _T_1392 = ~ _T_1390; // @[LZD.scala 49:27]
  assign _T_1393 = _T_1389 | _T_1392; // @[LZD.scala 49:25]
  assign _T_1394 = _T_1381[0:0]; // @[LZD.scala 49:47]
  assign _T_1395 = _T_1388[0:0]; // @[LZD.scala 49:59]
  assign _T_1396 = _T_1389 ? _T_1394 : _T_1395; // @[LZD.scala 49:35]
  assign _T_1398 = {_T_1391,_T_1393,_T_1396}; // @[Cat.scala 29:58]
  assign _T_1399 = _T_1373[2]; // @[Shift.scala 12:21]
  assign _T_1400 = _T_1398[2]; // @[Shift.scala 12:21]
  assign _T_1401 = _T_1399 | _T_1400; // @[LZD.scala 49:16]
  assign _T_1402 = ~ _T_1400; // @[LZD.scala 49:27]
  assign _T_1403 = _T_1399 | _T_1402; // @[LZD.scala 49:25]
  assign _T_1404 = _T_1373[1:0]; // @[LZD.scala 49:47]
  assign _T_1405 = _T_1398[1:0]; // @[LZD.scala 49:59]
  assign _T_1406 = _T_1399 ? _T_1404 : _T_1405; // @[LZD.scala 49:35]
  assign _T_1408 = {_T_1401,_T_1403,_T_1406}; // @[Cat.scala 29:58]
  assign _T_1409 = _T_1347[7:0]; // @[LZD.scala 44:32]
  assign _T_1410 = _T_1409[7:4]; // @[LZD.scala 43:32]
  assign _T_1411 = _T_1410[3:2]; // @[LZD.scala 43:32]
  assign _T_1412 = _T_1411 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1413 = _T_1411[1]; // @[LZD.scala 39:21]
  assign _T_1414 = _T_1411[0]; // @[LZD.scala 39:30]
  assign _T_1415 = ~ _T_1414; // @[LZD.scala 39:27]
  assign _T_1416 = _T_1413 | _T_1415; // @[LZD.scala 39:25]
  assign _T_1417 = {_T_1412,_T_1416}; // @[Cat.scala 29:58]
  assign _T_1418 = _T_1410[1:0]; // @[LZD.scala 44:32]
  assign _T_1419 = _T_1418 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1420 = _T_1418[1]; // @[LZD.scala 39:21]
  assign _T_1421 = _T_1418[0]; // @[LZD.scala 39:30]
  assign _T_1422 = ~ _T_1421; // @[LZD.scala 39:27]
  assign _T_1423 = _T_1420 | _T_1422; // @[LZD.scala 39:25]
  assign _T_1424 = {_T_1419,_T_1423}; // @[Cat.scala 29:58]
  assign _T_1425 = _T_1417[1]; // @[Shift.scala 12:21]
  assign _T_1426 = _T_1424[1]; // @[Shift.scala 12:21]
  assign _T_1427 = _T_1425 | _T_1426; // @[LZD.scala 49:16]
  assign _T_1428 = ~ _T_1426; // @[LZD.scala 49:27]
  assign _T_1429 = _T_1425 | _T_1428; // @[LZD.scala 49:25]
  assign _T_1430 = _T_1417[0:0]; // @[LZD.scala 49:47]
  assign _T_1431 = _T_1424[0:0]; // @[LZD.scala 49:59]
  assign _T_1432 = _T_1425 ? _T_1430 : _T_1431; // @[LZD.scala 49:35]
  assign _T_1434 = {_T_1427,_T_1429,_T_1432}; // @[Cat.scala 29:58]
  assign _T_1435 = _T_1409[3:0]; // @[LZD.scala 44:32]
  assign _T_1436 = _T_1435[3:2]; // @[LZD.scala 43:32]
  assign _T_1437 = _T_1436 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1438 = _T_1436[1]; // @[LZD.scala 39:21]
  assign _T_1439 = _T_1436[0]; // @[LZD.scala 39:30]
  assign _T_1440 = ~ _T_1439; // @[LZD.scala 39:27]
  assign _T_1441 = _T_1438 | _T_1440; // @[LZD.scala 39:25]
  assign _T_1442 = {_T_1437,_T_1441}; // @[Cat.scala 29:58]
  assign _T_1443 = _T_1435[1:0]; // @[LZD.scala 44:32]
  assign _T_1444 = _T_1443 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1445 = _T_1443[1]; // @[LZD.scala 39:21]
  assign _T_1446 = _T_1443[0]; // @[LZD.scala 39:30]
  assign _T_1447 = ~ _T_1446; // @[LZD.scala 39:27]
  assign _T_1448 = _T_1445 | _T_1447; // @[LZD.scala 39:25]
  assign _T_1449 = {_T_1444,_T_1448}; // @[Cat.scala 29:58]
  assign _T_1450 = _T_1442[1]; // @[Shift.scala 12:21]
  assign _T_1451 = _T_1449[1]; // @[Shift.scala 12:21]
  assign _T_1452 = _T_1450 | _T_1451; // @[LZD.scala 49:16]
  assign _T_1453 = ~ _T_1451; // @[LZD.scala 49:27]
  assign _T_1454 = _T_1450 | _T_1453; // @[LZD.scala 49:25]
  assign _T_1455 = _T_1442[0:0]; // @[LZD.scala 49:47]
  assign _T_1456 = _T_1449[0:0]; // @[LZD.scala 49:59]
  assign _T_1457 = _T_1450 ? _T_1455 : _T_1456; // @[LZD.scala 49:35]
  assign _T_1459 = {_T_1452,_T_1454,_T_1457}; // @[Cat.scala 29:58]
  assign _T_1460 = _T_1434[2]; // @[Shift.scala 12:21]
  assign _T_1461 = _T_1459[2]; // @[Shift.scala 12:21]
  assign _T_1462 = _T_1460 | _T_1461; // @[LZD.scala 49:16]
  assign _T_1463 = ~ _T_1461; // @[LZD.scala 49:27]
  assign _T_1464 = _T_1460 | _T_1463; // @[LZD.scala 49:25]
  assign _T_1465 = _T_1434[1:0]; // @[LZD.scala 49:47]
  assign _T_1466 = _T_1459[1:0]; // @[LZD.scala 49:59]
  assign _T_1467 = _T_1460 ? _T_1465 : _T_1466; // @[LZD.scala 49:35]
  assign _T_1469 = {_T_1462,_T_1464,_T_1467}; // @[Cat.scala 29:58]
  assign _T_1470 = _T_1408[3]; // @[Shift.scala 12:21]
  assign _T_1471 = _T_1469[3]; // @[Shift.scala 12:21]
  assign _T_1472 = _T_1470 | _T_1471; // @[LZD.scala 49:16]
  assign _T_1473 = ~ _T_1471; // @[LZD.scala 49:27]
  assign _T_1474 = _T_1470 | _T_1473; // @[LZD.scala 49:25]
  assign _T_1475 = _T_1408[2:0]; // @[LZD.scala 49:47]
  assign _T_1476 = _T_1469[2:0]; // @[LZD.scala 49:59]
  assign _T_1477 = _T_1470 ? _T_1475 : _T_1476; // @[LZD.scala 49:35]
  assign _T_1479 = {_T_1472,_T_1474,_T_1477}; // @[Cat.scala 29:58]
  assign _T_1480 = _T_1346[10:0]; // @[LZD.scala 44:32]
  assign _T_1481 = _T_1480[10:3]; // @[LZD.scala 43:32]
  assign _T_1482 = _T_1481[7:4]; // @[LZD.scala 43:32]
  assign _T_1483 = _T_1482[3:2]; // @[LZD.scala 43:32]
  assign _T_1484 = _T_1483 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1485 = _T_1483[1]; // @[LZD.scala 39:21]
  assign _T_1486 = _T_1483[0]; // @[LZD.scala 39:30]
  assign _T_1487 = ~ _T_1486; // @[LZD.scala 39:27]
  assign _T_1488 = _T_1485 | _T_1487; // @[LZD.scala 39:25]
  assign _T_1489 = {_T_1484,_T_1488}; // @[Cat.scala 29:58]
  assign _T_1490 = _T_1482[1:0]; // @[LZD.scala 44:32]
  assign _T_1491 = _T_1490 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1492 = _T_1490[1]; // @[LZD.scala 39:21]
  assign _T_1493 = _T_1490[0]; // @[LZD.scala 39:30]
  assign _T_1494 = ~ _T_1493; // @[LZD.scala 39:27]
  assign _T_1495 = _T_1492 | _T_1494; // @[LZD.scala 39:25]
  assign _T_1496 = {_T_1491,_T_1495}; // @[Cat.scala 29:58]
  assign _T_1497 = _T_1489[1]; // @[Shift.scala 12:21]
  assign _T_1498 = _T_1496[1]; // @[Shift.scala 12:21]
  assign _T_1499 = _T_1497 | _T_1498; // @[LZD.scala 49:16]
  assign _T_1500 = ~ _T_1498; // @[LZD.scala 49:27]
  assign _T_1501 = _T_1497 | _T_1500; // @[LZD.scala 49:25]
  assign _T_1502 = _T_1489[0:0]; // @[LZD.scala 49:47]
  assign _T_1503 = _T_1496[0:0]; // @[LZD.scala 49:59]
  assign _T_1504 = _T_1497 ? _T_1502 : _T_1503; // @[LZD.scala 49:35]
  assign _T_1506 = {_T_1499,_T_1501,_T_1504}; // @[Cat.scala 29:58]
  assign _T_1507 = _T_1481[3:0]; // @[LZD.scala 44:32]
  assign _T_1508 = _T_1507[3:2]; // @[LZD.scala 43:32]
  assign _T_1509 = _T_1508 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1510 = _T_1508[1]; // @[LZD.scala 39:21]
  assign _T_1511 = _T_1508[0]; // @[LZD.scala 39:30]
  assign _T_1512 = ~ _T_1511; // @[LZD.scala 39:27]
  assign _T_1513 = _T_1510 | _T_1512; // @[LZD.scala 39:25]
  assign _T_1514 = {_T_1509,_T_1513}; // @[Cat.scala 29:58]
  assign _T_1515 = _T_1507[1:0]; // @[LZD.scala 44:32]
  assign _T_1516 = _T_1515 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1517 = _T_1515[1]; // @[LZD.scala 39:21]
  assign _T_1518 = _T_1515[0]; // @[LZD.scala 39:30]
  assign _T_1519 = ~ _T_1518; // @[LZD.scala 39:27]
  assign _T_1520 = _T_1517 | _T_1519; // @[LZD.scala 39:25]
  assign _T_1521 = {_T_1516,_T_1520}; // @[Cat.scala 29:58]
  assign _T_1522 = _T_1514[1]; // @[Shift.scala 12:21]
  assign _T_1523 = _T_1521[1]; // @[Shift.scala 12:21]
  assign _T_1524 = _T_1522 | _T_1523; // @[LZD.scala 49:16]
  assign _T_1525 = ~ _T_1523; // @[LZD.scala 49:27]
  assign _T_1526 = _T_1522 | _T_1525; // @[LZD.scala 49:25]
  assign _T_1527 = _T_1514[0:0]; // @[LZD.scala 49:47]
  assign _T_1528 = _T_1521[0:0]; // @[LZD.scala 49:59]
  assign _T_1529 = _T_1522 ? _T_1527 : _T_1528; // @[LZD.scala 49:35]
  assign _T_1531 = {_T_1524,_T_1526,_T_1529}; // @[Cat.scala 29:58]
  assign _T_1532 = _T_1506[2]; // @[Shift.scala 12:21]
  assign _T_1533 = _T_1531[2]; // @[Shift.scala 12:21]
  assign _T_1534 = _T_1532 | _T_1533; // @[LZD.scala 49:16]
  assign _T_1535 = ~ _T_1533; // @[LZD.scala 49:27]
  assign _T_1536 = _T_1532 | _T_1535; // @[LZD.scala 49:25]
  assign _T_1537 = _T_1506[1:0]; // @[LZD.scala 49:47]
  assign _T_1538 = _T_1531[1:0]; // @[LZD.scala 49:59]
  assign _T_1539 = _T_1532 ? _T_1537 : _T_1538; // @[LZD.scala 49:35]
  assign _T_1541 = {_T_1534,_T_1536,_T_1539}; // @[Cat.scala 29:58]
  assign _T_1542 = _T_1480[2:0]; // @[LZD.scala 44:32]
  assign _T_1543 = _T_1542[2:1]; // @[LZD.scala 43:32]
  assign _T_1544 = _T_1543 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1545 = _T_1543[1]; // @[LZD.scala 39:21]
  assign _T_1546 = _T_1543[0]; // @[LZD.scala 39:30]
  assign _T_1547 = ~ _T_1546; // @[LZD.scala 39:27]
  assign _T_1548 = _T_1545 | _T_1547; // @[LZD.scala 39:25]
  assign _T_1549 = {_T_1544,_T_1548}; // @[Cat.scala 29:58]
  assign _T_1550 = _T_1542[0:0]; // @[LZD.scala 44:32]
  assign _T_1552 = _T_1549[1]; // @[Shift.scala 12:21]
  assign _T_1554 = _T_1549[0:0]; // @[LZD.scala 55:32]
  assign _T_1555 = _T_1552 ? _T_1554 : _T_1550; // @[LZD.scala 55:20]
  assign _T_1557 = _T_1541[3]; // @[Shift.scala 12:21]
  assign _T_1559 = {1'h1,_T_1552,_T_1555}; // @[Cat.scala 29:58]
  assign _T_1560 = _T_1541[2:0]; // @[LZD.scala 55:32]
  assign _T_1561 = _T_1557 ? _T_1560 : _T_1559; // @[LZD.scala 55:20]
  assign _T_1562 = {_T_1557,_T_1561}; // @[Cat.scala 29:58]
  assign _T_1563 = _T_1479[4]; // @[Shift.scala 12:21]
  assign _T_1565 = _T_1479[3:0]; // @[LZD.scala 55:32]
  assign _T_1566 = _T_1563 ? _T_1565 : _T_1562; // @[LZD.scala 55:20]
  assign _T_1567 = {_T_1563,_T_1566}; // @[Cat.scala 29:58]
  assign _T_1568 = _T_1345[5]; // @[Shift.scala 12:21]
  assign _T_1570 = _T_1345[4:0]; // @[LZD.scala 55:32]
  assign _T_1571 = _T_1568 ? _T_1570 : _T_1567; // @[LZD.scala 55:20]
  assign sumLZD = {_T_1568,_T_1571}; // @[Cat.scala 29:58]
  assign shiftValue = ~ sumLZD; // @[PositFMA.scala 126:24]
  assign _T_1572 = signSumSig[57:0]; // @[PositFMA.scala 127:38]
  assign _T_1573 = shiftValue < 6'h3a; // @[Shift.scala 16:24]
  assign _T_1575 = shiftValue[5]; // @[Shift.scala 12:21]
  assign _T_1576 = _T_1572[25:0]; // @[Shift.scala 64:52]
  assign _T_1578 = {_T_1576,32'h0}; // @[Cat.scala 29:58]
  assign _T_1579 = _T_1575 ? _T_1578 : _T_1572; // @[Shift.scala 64:27]
  assign _T_1580 = shiftValue[4:0]; // @[Shift.scala 66:70]
  assign _T_1581 = _T_1580[4]; // @[Shift.scala 12:21]
  assign _T_1582 = _T_1579[41:0]; // @[Shift.scala 64:52]
  assign _T_1584 = {_T_1582,16'h0}; // @[Cat.scala 29:58]
  assign _T_1585 = _T_1581 ? _T_1584 : _T_1579; // @[Shift.scala 64:27]
  assign _T_1586 = _T_1580[3:0]; // @[Shift.scala 66:70]
  assign _T_1587 = _T_1586[3]; // @[Shift.scala 12:21]
  assign _T_1588 = _T_1585[49:0]; // @[Shift.scala 64:52]
  assign _T_1590 = {_T_1588,8'h0}; // @[Cat.scala 29:58]
  assign _T_1591 = _T_1587 ? _T_1590 : _T_1585; // @[Shift.scala 64:27]
  assign _T_1592 = _T_1586[2:0]; // @[Shift.scala 66:70]
  assign _T_1593 = _T_1592[2]; // @[Shift.scala 12:21]
  assign _T_1594 = _T_1591[53:0]; // @[Shift.scala 64:52]
  assign _T_1596 = {_T_1594,4'h0}; // @[Cat.scala 29:58]
  assign _T_1597 = _T_1593 ? _T_1596 : _T_1591; // @[Shift.scala 64:27]
  assign _T_1598 = _T_1592[1:0]; // @[Shift.scala 66:70]
  assign _T_1599 = _T_1598[1]; // @[Shift.scala 12:21]
  assign _T_1600 = _T_1597[55:0]; // @[Shift.scala 64:52]
  assign _T_1602 = {_T_1600,2'h0}; // @[Cat.scala 29:58]
  assign _T_1603 = _T_1599 ? _T_1602 : _T_1597; // @[Shift.scala 64:27]
  assign _T_1604 = _T_1598[0:0]; // @[Shift.scala 66:70]
  assign _T_1606 = _T_1603[56:0]; // @[Shift.scala 64:52]
  assign _T_1607 = {_T_1606,1'h0}; // @[Cat.scala 29:58]
  assign _T_1608 = _T_1604 ? _T_1607 : _T_1603; // @[Shift.scala 64:27]
  assign normalFracTmp = _T_1573 ? _T_1608 : 58'h0; // @[Shift.scala 16:10]
  assign _T_1610 = $signed(greaterScale) + $signed(8'sh2); // @[PositFMA.scala 130:36]
  assign _T_1611 = $signed(_T_1610); // @[PositFMA.scala 130:36]
  assign _T_1612 = {1'h1,_T_1568,_T_1571}; // @[Cat.scala 29:58]
  assign _T_1613 = $signed(_T_1612); // @[PositFMA.scala 130:61]
  assign _GEN_20 = {{1{_T_1613[6]}},_T_1613}; // @[PositFMA.scala 130:42]
  assign _T_1615 = $signed(_T_1611) + $signed(_GEN_20); // @[PositFMA.scala 130:42]
  assign sumScale = $signed(_T_1615); // @[PositFMA.scala 130:42]
  assign sumFrac = normalFracTmp[57:30]; // @[PositFMA.scala 131:41]
  assign grsTmp = normalFracTmp[29:0]; // @[PositFMA.scala 134:41]
  assign _T_1616 = grsTmp[29:28]; // @[PositFMA.scala 137:40]
  assign _T_1617 = grsTmp[27:0]; // @[PositFMA.scala 137:56]
  assign _T_1618 = _T_1617 != 28'h0; // @[PositFMA.scala 137:60]
  assign underflow = $signed(sumScale) < $signed(-8'sh3d); // @[PositFMA.scala 144:32]
  assign overflow = $signed(sumScale) > $signed(8'sh3c); // @[PositFMA.scala 145:32]
  assign _T_1619 = signSumSig != 60'h0; // @[PositFMA.scala 154:32]
  assign decF_isZero = ~ _T_1619; // @[PositFMA.scala 154:20]
  assign _T_1621 = underflow ? $signed(-8'sh3d) : $signed(sumScale); // @[Mux.scala 87:16]
  assign _T_1622 = overflow ? $signed(8'sh3c) : $signed(_T_1621); // @[Mux.scala 87:16]
  assign _GEN_21 = _T_1622[6:0]; // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  assign decF_scale = $signed(_GEN_21); // @[PositFMA.scala 151:18 PositFMA.scala 157:17]
  assign _T_1623 = decF_scale[0]; // @[convert.scala 46:61]
  assign _T_1624 = ~ _T_1623; // @[convert.scala 46:52]
  assign _T_1626 = sumSign ? _T_1624 : _T_1623; // @[convert.scala 46:42]
  assign _T_1627 = decF_scale[6:1]; // @[convert.scala 48:34]
  assign _T_1628 = _T_1627[5:5]; // @[convert.scala 49:36]
  assign _T_1630 = ~ _T_1627; // @[convert.scala 50:36]
  assign _T_1631 = $signed(_T_1630); // @[convert.scala 50:36]
  assign _T_1632 = _T_1628 ? $signed(_T_1631) : $signed(_T_1627); // @[convert.scala 50:28]
  assign _T_1633 = _T_1628 ^ sumSign; // @[convert.scala 51:31]
  assign _T_1634 = ~ _T_1633; // @[convert.scala 52:43]
  assign _T_1638 = {_T_1634,_T_1633,_T_1626,sumFrac,_T_1616,_T_1618}; // @[Cat.scala 29:58]
  assign _T_1639 = $unsigned(_T_1632); // @[Shift.scala 39:17]
  assign _T_1640 = _T_1639 < 6'h22; // @[Shift.scala 39:24]
  assign _T_1642 = _T_1638[33:32]; // @[Shift.scala 90:30]
  assign _T_1643 = _T_1638[31:0]; // @[Shift.scala 90:48]
  assign _T_1644 = _T_1643 != 32'h0; // @[Shift.scala 90:57]
  assign _GEN_22 = {{1'd0}, _T_1644}; // @[Shift.scala 90:39]
  assign _T_1645 = _T_1642 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_1646 = _T_1639[5]; // @[Shift.scala 12:21]
  assign _T_1647 = _T_1638[33]; // @[Shift.scala 12:21]
  assign _T_1649 = _T_1647 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 71:12]
  assign _T_1650 = {_T_1649,_T_1645}; // @[Cat.scala 29:58]
  assign _T_1651 = _T_1646 ? _T_1650 : _T_1638; // @[Shift.scala 91:22]
  assign _T_1652 = _T_1639[4:0]; // @[Shift.scala 92:77]
  assign _T_1653 = _T_1651[33:16]; // @[Shift.scala 90:30]
  assign _T_1654 = _T_1651[15:0]; // @[Shift.scala 90:48]
  assign _T_1655 = _T_1654 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_23 = {{17'd0}, _T_1655}; // @[Shift.scala 90:39]
  assign _T_1656 = _T_1653 | _GEN_23; // @[Shift.scala 90:39]
  assign _T_1657 = _T_1652[4]; // @[Shift.scala 12:21]
  assign _T_1658 = _T_1651[33]; // @[Shift.scala 12:21]
  assign _T_1660 = _T_1658 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_1661 = {_T_1660,_T_1656}; // @[Cat.scala 29:58]
  assign _T_1662 = _T_1657 ? _T_1661 : _T_1651; // @[Shift.scala 91:22]
  assign _T_1663 = _T_1652[3:0]; // @[Shift.scala 92:77]
  assign _T_1664 = _T_1662[33:8]; // @[Shift.scala 90:30]
  assign _T_1665 = _T_1662[7:0]; // @[Shift.scala 90:48]
  assign _T_1666 = _T_1665 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_24 = {{25'd0}, _T_1666}; // @[Shift.scala 90:39]
  assign _T_1667 = _T_1664 | _GEN_24; // @[Shift.scala 90:39]
  assign _T_1668 = _T_1663[3]; // @[Shift.scala 12:21]
  assign _T_1669 = _T_1662[33]; // @[Shift.scala 12:21]
  assign _T_1671 = _T_1669 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_1672 = {_T_1671,_T_1667}; // @[Cat.scala 29:58]
  assign _T_1673 = _T_1668 ? _T_1672 : _T_1662; // @[Shift.scala 91:22]
  assign _T_1674 = _T_1663[2:0]; // @[Shift.scala 92:77]
  assign _T_1675 = _T_1673[33:4]; // @[Shift.scala 90:30]
  assign _T_1676 = _T_1673[3:0]; // @[Shift.scala 90:48]
  assign _T_1677 = _T_1676 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_25 = {{29'd0}, _T_1677}; // @[Shift.scala 90:39]
  assign _T_1678 = _T_1675 | _GEN_25; // @[Shift.scala 90:39]
  assign _T_1679 = _T_1674[2]; // @[Shift.scala 12:21]
  assign _T_1680 = _T_1673[33]; // @[Shift.scala 12:21]
  assign _T_1682 = _T_1680 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_1683 = {_T_1682,_T_1678}; // @[Cat.scala 29:58]
  assign _T_1684 = _T_1679 ? _T_1683 : _T_1673; // @[Shift.scala 91:22]
  assign _T_1685 = _T_1674[1:0]; // @[Shift.scala 92:77]
  assign _T_1686 = _T_1684[33:2]; // @[Shift.scala 90:30]
  assign _T_1687 = _T_1684[1:0]; // @[Shift.scala 90:48]
  assign _T_1688 = _T_1687 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_26 = {{31'd0}, _T_1688}; // @[Shift.scala 90:39]
  assign _T_1689 = _T_1686 | _GEN_26; // @[Shift.scala 90:39]
  assign _T_1690 = _T_1685[1]; // @[Shift.scala 12:21]
  assign _T_1691 = _T_1684[33]; // @[Shift.scala 12:21]
  assign _T_1693 = _T_1691 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_1694 = {_T_1693,_T_1689}; // @[Cat.scala 29:58]
  assign _T_1695 = _T_1690 ? _T_1694 : _T_1684; // @[Shift.scala 91:22]
  assign _T_1696 = _T_1685[0:0]; // @[Shift.scala 92:77]
  assign _T_1697 = _T_1695[33:1]; // @[Shift.scala 90:30]
  assign _T_1698 = _T_1695[0:0]; // @[Shift.scala 90:48]
  assign _GEN_27 = {{32'd0}, _T_1698}; // @[Shift.scala 90:39]
  assign _T_1700 = _T_1697 | _GEN_27; // @[Shift.scala 90:39]
  assign _T_1702 = _T_1695[33]; // @[Shift.scala 12:21]
  assign _T_1703 = {_T_1702,_T_1700}; // @[Cat.scala 29:58]
  assign _T_1704 = _T_1696 ? _T_1703 : _T_1695; // @[Shift.scala 91:22]
  assign _T_1707 = _T_1647 ? 34'h3ffffffff : 34'h0; // @[Bitwise.scala 71:12]
  assign _T_1708 = _T_1640 ? _T_1704 : _T_1707; // @[Shift.scala 39:10]
  assign _T_1709 = _T_1708[3]; // @[convert.scala 55:31]
  assign _T_1710 = _T_1708[2]; // @[convert.scala 56:31]
  assign _T_1711 = _T_1708[1]; // @[convert.scala 57:31]
  assign _T_1712 = _T_1708[0]; // @[convert.scala 58:31]
  assign _T_1713 = _T_1708[33:3]; // @[convert.scala 59:69]
  assign _T_1714 = _T_1713 != 31'h0; // @[convert.scala 59:81]
  assign _T_1715 = ~ _T_1714; // @[convert.scala 59:50]
  assign _T_1717 = _T_1713 == 31'h7fffffff; // @[convert.scala 60:81]
  assign _T_1718 = _T_1709 | _T_1711; // @[convert.scala 61:44]
  assign _T_1719 = _T_1718 | _T_1712; // @[convert.scala 61:52]
  assign _T_1720 = _T_1710 & _T_1719; // @[convert.scala 61:36]
  assign _T_1721 = ~ _T_1717; // @[convert.scala 62:63]
  assign _T_1722 = _T_1721 & _T_1720; // @[convert.scala 62:103]
  assign _T_1723 = _T_1715 | _T_1722; // @[convert.scala 62:60]
  assign _GEN_28 = {{30'd0}, _T_1723}; // @[convert.scala 63:56]
  assign _T_1726 = _T_1713 + _GEN_28; // @[convert.scala 63:56]
  assign _T_1727 = {sumSign,_T_1726}; // @[Cat.scala 29:58]
  assign io_F = _T_1735; // @[PositFMA.scala 174:15]
  assign io_outValid = _T_1731; // @[PositFMA.scala 173:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  outIsNaR_phase2 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  mulSig_phase2 = _RAND_1[58:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  addFrac_phase2 = _RAND_2[27:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mulScale_phase2 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addScale_phase2 = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addSign_phase2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addZero_phase2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  inValid_phase2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1731 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_1735 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (io_inValid) begin
      outIsNaR_phase2 <= outIsNaR;
    end
    if (io_inValid) begin
      mulSig_phase2 <= mulSig;
    end
    if (io_inValid) begin
      addFrac_phase2 <= decC_fraction;
    end
    if (io_inValid) begin
      mulScale_phase2 <= mulScale;
    end
    if (io_inValid) begin
      addScale_phase2 <= decC_scale;
    end
    if (io_inValid) begin
      addSign_phase2 <= _T_627;
    end
    if (io_inValid) begin
      addZero_phase2 <= decC_isZero;
    end
    if (reset) begin
      inValid_phase2 <= 1'h0;
    end else begin
      inValid_phase2 <= io_inValid;
    end
    if (reset) begin
      _T_1731 <= 1'h0;
    end else begin
      _T_1731 <= inValid_phase2;
    end
    if (inValid_phase2) begin
      if (outIsNaR_phase2) begin
        _T_1735 <= 32'h80000000;
      end else begin
        if (decF_isZero) begin
          _T_1735 <= 32'h0;
        end else begin
          _T_1735 <= _T_1727;
        end
      end
    end
  end
endmodule
