module PositAdder8_1(
  input        clock,
  input        reset,
  input  [7:0] io_A,
  input  [7:0] io_B,
  output [7:0] io_S
);
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [5:0] _T_4; // @[convert.scala 19:24]
  wire [5:0] _T_5; // @[convert.scala 19:43]
  wire [5:0] _T_6; // @[convert.scala 19:39]
  wire [3:0] _T_7; // @[LZD.scala 43:32]
  wire [1:0] _T_8; // @[LZD.scala 43:32]
  wire  _T_9; // @[LZD.scala 39:14]
  wire  _T_10; // @[LZD.scala 39:21]
  wire  _T_11; // @[LZD.scala 39:30]
  wire  _T_12; // @[LZD.scala 39:27]
  wire  _T_13; // @[LZD.scala 39:25]
  wire [1:0] _T_14; // @[Cat.scala 29:58]
  wire [1:0] _T_15; // @[LZD.scala 44:32]
  wire  _T_16; // @[LZD.scala 39:14]
  wire  _T_17; // @[LZD.scala 39:21]
  wire  _T_18; // @[LZD.scala 39:30]
  wire  _T_19; // @[LZD.scala 39:27]
  wire  _T_20; // @[LZD.scala 39:25]
  wire [1:0] _T_21; // @[Cat.scala 29:58]
  wire  _T_22; // @[Shift.scala 12:21]
  wire  _T_23; // @[Shift.scala 12:21]
  wire  _T_24; // @[LZD.scala 49:16]
  wire  _T_25; // @[LZD.scala 49:27]
  wire  _T_26; // @[LZD.scala 49:25]
  wire  _T_27; // @[LZD.scala 49:47]
  wire  _T_28; // @[LZD.scala 49:59]
  wire  _T_29; // @[LZD.scala 49:35]
  wire [2:0] _T_31; // @[Cat.scala 29:58]
  wire [1:0] _T_32; // @[LZD.scala 44:32]
  wire  _T_33; // @[LZD.scala 39:14]
  wire  _T_34; // @[LZD.scala 39:21]
  wire  _T_35; // @[LZD.scala 39:30]
  wire  _T_36; // @[LZD.scala 39:27]
  wire  _T_37; // @[LZD.scala 39:25]
  wire [1:0] _T_38; // @[Cat.scala 29:58]
  wire  _T_39; // @[Shift.scala 12:21]
  wire [1:0] _T_41; // @[LZD.scala 55:32]
  wire [1:0] _T_42; // @[LZD.scala 55:20]
  wire [2:0] _T_43; // @[Cat.scala 29:58]
  wire [2:0] _T_44; // @[convert.scala 21:22]
  wire [4:0] _T_45; // @[convert.scala 22:36]
  wire  _T_46; // @[Shift.scala 16:24]
  wire  _T_48; // @[Shift.scala 12:21]
  wire  _T_49; // @[Shift.scala 64:52]
  wire [4:0] _T_51; // @[Cat.scala 29:58]
  wire [4:0] _T_52; // @[Shift.scala 64:27]
  wire [1:0] _T_53; // @[Shift.scala 66:70]
  wire  _T_54; // @[Shift.scala 12:21]
  wire [2:0] _T_55; // @[Shift.scala 64:52]
  wire [4:0] _T_57; // @[Cat.scala 29:58]
  wire [4:0] _T_58; // @[Shift.scala 64:27]
  wire  _T_59; // @[Shift.scala 66:70]
  wire [3:0] _T_61; // @[Shift.scala 64:52]
  wire [4:0] _T_62; // @[Cat.scala 29:58]
  wire [4:0] _T_63; // @[Shift.scala 64:27]
  wire [4:0] _T_64; // @[Shift.scala 16:10]
  wire  _T_65; // @[convert.scala 23:34]
  wire [3:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_67; // @[convert.scala 25:26]
  wire [2:0] _T_69; // @[convert.scala 25:42]
  wire  _T_72; // @[convert.scala 26:67]
  wire  _T_73; // @[convert.scala 26:51]
  wire [4:0] _T_74; // @[Cat.scala 29:58]
  wire [6:0] _T_76; // @[convert.scala 29:56]
  wire  _T_77; // @[convert.scala 29:60]
  wire  _T_78; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_81; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [4:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_90; // @[convert.scala 18:24]
  wire  _T_91; // @[convert.scala 18:40]
  wire  _T_92; // @[convert.scala 18:36]
  wire [5:0] _T_93; // @[convert.scala 19:24]
  wire [5:0] _T_94; // @[convert.scala 19:43]
  wire [5:0] _T_95; // @[convert.scala 19:39]
  wire [3:0] _T_96; // @[LZD.scala 43:32]
  wire [1:0] _T_97; // @[LZD.scala 43:32]
  wire  _T_98; // @[LZD.scala 39:14]
  wire  _T_99; // @[LZD.scala 39:21]
  wire  _T_100; // @[LZD.scala 39:30]
  wire  _T_101; // @[LZD.scala 39:27]
  wire  _T_102; // @[LZD.scala 39:25]
  wire [1:0] _T_103; // @[Cat.scala 29:58]
  wire [1:0] _T_104; // @[LZD.scala 44:32]
  wire  _T_105; // @[LZD.scala 39:14]
  wire  _T_106; // @[LZD.scala 39:21]
  wire  _T_107; // @[LZD.scala 39:30]
  wire  _T_108; // @[LZD.scala 39:27]
  wire  _T_109; // @[LZD.scala 39:25]
  wire [1:0] _T_110; // @[Cat.scala 29:58]
  wire  _T_111; // @[Shift.scala 12:21]
  wire  _T_112; // @[Shift.scala 12:21]
  wire  _T_113; // @[LZD.scala 49:16]
  wire  _T_114; // @[LZD.scala 49:27]
  wire  _T_115; // @[LZD.scala 49:25]
  wire  _T_116; // @[LZD.scala 49:47]
  wire  _T_117; // @[LZD.scala 49:59]
  wire  _T_118; // @[LZD.scala 49:35]
  wire [2:0] _T_120; // @[Cat.scala 29:58]
  wire [1:0] _T_121; // @[LZD.scala 44:32]
  wire  _T_122; // @[LZD.scala 39:14]
  wire  _T_123; // @[LZD.scala 39:21]
  wire  _T_124; // @[LZD.scala 39:30]
  wire  _T_125; // @[LZD.scala 39:27]
  wire  _T_126; // @[LZD.scala 39:25]
  wire [1:0] _T_127; // @[Cat.scala 29:58]
  wire  _T_128; // @[Shift.scala 12:21]
  wire [1:0] _T_130; // @[LZD.scala 55:32]
  wire [1:0] _T_131; // @[LZD.scala 55:20]
  wire [2:0] _T_132; // @[Cat.scala 29:58]
  wire [2:0] _T_133; // @[convert.scala 21:22]
  wire [4:0] _T_134; // @[convert.scala 22:36]
  wire  _T_135; // @[Shift.scala 16:24]
  wire  _T_137; // @[Shift.scala 12:21]
  wire  _T_138; // @[Shift.scala 64:52]
  wire [4:0] _T_140; // @[Cat.scala 29:58]
  wire [4:0] _T_141; // @[Shift.scala 64:27]
  wire [1:0] _T_142; // @[Shift.scala 66:70]
  wire  _T_143; // @[Shift.scala 12:21]
  wire [2:0] _T_144; // @[Shift.scala 64:52]
  wire [4:0] _T_146; // @[Cat.scala 29:58]
  wire [4:0] _T_147; // @[Shift.scala 64:27]
  wire  _T_148; // @[Shift.scala 66:70]
  wire [3:0] _T_150; // @[Shift.scala 64:52]
  wire [4:0] _T_151; // @[Cat.scala 29:58]
  wire [4:0] _T_152; // @[Shift.scala 64:27]
  wire [4:0] _T_153; // @[Shift.scala 16:10]
  wire  _T_154; // @[convert.scala 23:34]
  wire [3:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_156; // @[convert.scala 25:26]
  wire [2:0] _T_158; // @[convert.scala 25:42]
  wire  _T_161; // @[convert.scala 26:67]
  wire  _T_162; // @[convert.scala 26:51]
  wire [4:0] _T_163; // @[Cat.scala 29:58]
  wire [6:0] _T_165; // @[convert.scala 29:56]
  wire  _T_166; // @[convert.scala 29:60]
  wire  _T_167; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_170; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [4:0] decB_scale; // @[convert.scala 32:24]
  wire  aGTb; // @[PositAdder.scala 24:32]
  wire  greaterSign; // @[PositAdder.scala 25:24]
  wire  smallerSign; // @[PositAdder.scala 26:24]
  wire [4:0] greaterExp; // @[PositAdder.scala 27:24]
  wire [4:0] smallerExp; // @[PositAdder.scala 28:24]
  wire [3:0] greaterFrac; // @[PositAdder.scala 29:24]
  wire [3:0] smallerFrac; // @[PositAdder.scala 30:24]
  wire  smallerZero; // @[PositAdder.scala 31:24]
  wire [4:0] _T_179; // @[PositAdder.scala 32:32]
  wire [4:0] scale_diff; // @[PositAdder.scala 32:32]
  wire  _T_180; // @[PositAdder.scala 33:38]
  wire [5:0] greaterSig; // @[Cat.scala 29:58]
  wire  _T_182; // @[PositAdder.scala 34:52]
  wire  _T_183; // @[PositAdder.scala 34:38]
  wire [8:0] _T_186; // @[Cat.scala 29:58]
  wire [4:0] _T_187; // @[PositAdder.scala 35:68]
  wire  _T_188; // @[Shift.scala 39:24]
  wire [3:0] _T_189; // @[Shift.scala 40:44]
  wire  _T_190; // @[Shift.scala 90:30]
  wire [7:0] _T_191; // @[Shift.scala 90:48]
  wire  _T_192; // @[Shift.scala 90:57]
  wire  _T_193; // @[Shift.scala 90:39]
  wire  _T_194; // @[Shift.scala 12:21]
  wire  _T_195; // @[Shift.scala 12:21]
  wire [7:0] _T_197; // @[Bitwise.scala 71:12]
  wire [8:0] _T_198; // @[Cat.scala 29:58]
  wire [8:0] _T_199; // @[Shift.scala 91:22]
  wire [2:0] _T_200; // @[Shift.scala 92:77]
  wire [4:0] _T_201; // @[Shift.scala 90:30]
  wire [3:0] _T_202; // @[Shift.scala 90:48]
  wire  _T_203; // @[Shift.scala 90:57]
  wire [4:0] _GEN_0; // @[Shift.scala 90:39]
  wire [4:0] _T_204; // @[Shift.scala 90:39]
  wire  _T_205; // @[Shift.scala 12:21]
  wire  _T_206; // @[Shift.scala 12:21]
  wire [3:0] _T_208; // @[Bitwise.scala 71:12]
  wire [8:0] _T_209; // @[Cat.scala 29:58]
  wire [8:0] _T_210; // @[Shift.scala 91:22]
  wire [1:0] _T_211; // @[Shift.scala 92:77]
  wire [6:0] _T_212; // @[Shift.scala 90:30]
  wire [1:0] _T_213; // @[Shift.scala 90:48]
  wire  _T_214; // @[Shift.scala 90:57]
  wire [6:0] _GEN_1; // @[Shift.scala 90:39]
  wire [6:0] _T_215; // @[Shift.scala 90:39]
  wire  _T_216; // @[Shift.scala 12:21]
  wire  _T_217; // @[Shift.scala 12:21]
  wire [1:0] _T_219; // @[Bitwise.scala 71:12]
  wire [8:0] _T_220; // @[Cat.scala 29:58]
  wire [8:0] _T_221; // @[Shift.scala 91:22]
  wire  _T_222; // @[Shift.scala 92:77]
  wire [7:0] _T_223; // @[Shift.scala 90:30]
  wire  _T_224; // @[Shift.scala 90:48]
  wire [7:0] _GEN_2; // @[Shift.scala 90:39]
  wire [7:0] _T_226; // @[Shift.scala 90:39]
  wire  _T_228; // @[Shift.scala 12:21]
  wire [8:0] _T_229; // @[Cat.scala 29:58]
  wire [8:0] _T_230; // @[Shift.scala 91:22]
  wire [8:0] _T_233; // @[Bitwise.scala 71:12]
  wire [8:0] smallerSig; // @[Shift.scala 39:10]
  wire [5:0] _T_234; // @[PositAdder.scala 36:45]
  wire [6:0] rawSumSig; // @[PositAdder.scala 36:32]
  wire  _T_235; // @[PositAdder.scala 37:31]
  wire  _T_236; // @[PositAdder.scala 37:59]
  wire  sumSign; // @[PositAdder.scala 37:43]
  wire [5:0] _T_237; // @[PositAdder.scala 38:48]
  wire [2:0] _T_238; // @[PositAdder.scala 38:63]
  wire [9:0] signSumSig; // @[Cat.scala 29:58]
  wire [8:0] _T_240; // @[PositAdder.scala 40:31]
  wire [8:0] _T_241; // @[PositAdder.scala 40:66]
  wire [8:0] sumXor; // @[PositAdder.scala 40:49]
  wire [7:0] _T_242; // @[LZD.scala 43:32]
  wire [3:0] _T_243; // @[LZD.scala 43:32]
  wire [1:0] _T_244; // @[LZD.scala 43:32]
  wire  _T_245; // @[LZD.scala 39:14]
  wire  _T_246; // @[LZD.scala 39:21]
  wire  _T_247; // @[LZD.scala 39:30]
  wire  _T_248; // @[LZD.scala 39:27]
  wire  _T_249; // @[LZD.scala 39:25]
  wire [1:0] _T_250; // @[Cat.scala 29:58]
  wire [1:0] _T_251; // @[LZD.scala 44:32]
  wire  _T_252; // @[LZD.scala 39:14]
  wire  _T_253; // @[LZD.scala 39:21]
  wire  _T_254; // @[LZD.scala 39:30]
  wire  _T_255; // @[LZD.scala 39:27]
  wire  _T_256; // @[LZD.scala 39:25]
  wire [1:0] _T_257; // @[Cat.scala 29:58]
  wire  _T_258; // @[Shift.scala 12:21]
  wire  _T_259; // @[Shift.scala 12:21]
  wire  _T_260; // @[LZD.scala 49:16]
  wire  _T_261; // @[LZD.scala 49:27]
  wire  _T_262; // @[LZD.scala 49:25]
  wire  _T_263; // @[LZD.scala 49:47]
  wire  _T_264; // @[LZD.scala 49:59]
  wire  _T_265; // @[LZD.scala 49:35]
  wire [2:0] _T_267; // @[Cat.scala 29:58]
  wire [3:0] _T_268; // @[LZD.scala 44:32]
  wire [1:0] _T_269; // @[LZD.scala 43:32]
  wire  _T_270; // @[LZD.scala 39:14]
  wire  _T_271; // @[LZD.scala 39:21]
  wire  _T_272; // @[LZD.scala 39:30]
  wire  _T_273; // @[LZD.scala 39:27]
  wire  _T_274; // @[LZD.scala 39:25]
  wire [1:0] _T_275; // @[Cat.scala 29:58]
  wire [1:0] _T_276; // @[LZD.scala 44:32]
  wire  _T_277; // @[LZD.scala 39:14]
  wire  _T_278; // @[LZD.scala 39:21]
  wire  _T_279; // @[LZD.scala 39:30]
  wire  _T_280; // @[LZD.scala 39:27]
  wire  _T_281; // @[LZD.scala 39:25]
  wire [1:0] _T_282; // @[Cat.scala 29:58]
  wire  _T_283; // @[Shift.scala 12:21]
  wire  _T_284; // @[Shift.scala 12:21]
  wire  _T_285; // @[LZD.scala 49:16]
  wire  _T_286; // @[LZD.scala 49:27]
  wire  _T_287; // @[LZD.scala 49:25]
  wire  _T_288; // @[LZD.scala 49:47]
  wire  _T_289; // @[LZD.scala 49:59]
  wire  _T_290; // @[LZD.scala 49:35]
  wire [2:0] _T_292; // @[Cat.scala 29:58]
  wire  _T_293; // @[Shift.scala 12:21]
  wire  _T_294; // @[Shift.scala 12:21]
  wire  _T_295; // @[LZD.scala 49:16]
  wire  _T_296; // @[LZD.scala 49:27]
  wire  _T_297; // @[LZD.scala 49:25]
  wire [1:0] _T_298; // @[LZD.scala 49:47]
  wire [1:0] _T_299; // @[LZD.scala 49:59]
  wire [1:0] _T_300; // @[LZD.scala 49:35]
  wire [3:0] _T_302; // @[Cat.scala 29:58]
  wire  _T_303; // @[LZD.scala 44:32]
  wire  _T_305; // @[Shift.scala 12:21]
  wire [2:0] _T_308; // @[Cat.scala 29:58]
  wire [2:0] _T_309; // @[LZD.scala 55:32]
  wire [2:0] _T_310; // @[LZD.scala 55:20]
  wire [3:0] sumLZD; // @[Cat.scala 29:58]
  wire [4:0] _T_311; // @[Cat.scala 29:58]
  wire [4:0] _T_312; // @[PositAdder.scala 42:38]
  wire [4:0] _T_314; // @[PositAdder.scala 42:45]
  wire [4:0] scaleBias; // @[PositAdder.scala 42:45]
  wire [5:0] sumScale; // @[PositAdder.scala 43:32]
  wire  overflow; // @[PositAdder.scala 44:30]
  wire [3:0] normalShift; // @[PositAdder.scala 45:22]
  wire [7:0] _T_315; // @[PositAdder.scala 46:36]
  wire  _T_316; // @[Shift.scala 16:24]
  wire [2:0] _T_317; // @[Shift.scala 17:37]
  wire  _T_318; // @[Shift.scala 12:21]
  wire [3:0] _T_319; // @[Shift.scala 64:52]
  wire [7:0] _T_321; // @[Cat.scala 29:58]
  wire [7:0] _T_322; // @[Shift.scala 64:27]
  wire [1:0] _T_323; // @[Shift.scala 66:70]
  wire  _T_324; // @[Shift.scala 12:21]
  wire [5:0] _T_325; // @[Shift.scala 64:52]
  wire [7:0] _T_327; // @[Cat.scala 29:58]
  wire [7:0] _T_328; // @[Shift.scala 64:27]
  wire  _T_329; // @[Shift.scala 66:70]
  wire [6:0] _T_331; // @[Shift.scala 64:52]
  wire [7:0] _T_332; // @[Cat.scala 29:58]
  wire [7:0] _T_333; // @[Shift.scala 64:27]
  wire [7:0] shiftSig; // @[Shift.scala 16:10]
  wire [5:0] _T_334; // @[PositAdder.scala 51:24]
  wire [3:0] decS_fraction; // @[PositAdder.scala 52:34]
  wire  decS_isNaR; // @[PositAdder.scala 53:32]
  wire  _T_337; // @[PositAdder.scala 54:33]
  wire  _T_338; // @[PositAdder.scala 54:21]
  wire  _T_339; // @[PositAdder.scala 54:52]
  wire  decS_isZero; // @[PositAdder.scala 54:37]
  wire [1:0] _T_341; // @[PositAdder.scala 55:33]
  wire  _T_342; // @[PositAdder.scala 55:49]
  wire  _T_343; // @[PositAdder.scala 55:63]
  wire  _T_344; // @[PositAdder.scala 55:53]
  wire [4:0] _GEN_3; // @[PositAdder.scala 48:25 PositAdder.scala 51:18]
  wire [4:0] decS_scale; // @[PositAdder.scala 48:25 PositAdder.scala 51:18]
  wire  _T_347; // @[convert.scala 46:61]
  wire  _T_348; // @[convert.scala 46:52]
  wire  _T_350; // @[convert.scala 46:42]
  wire [3:0] _T_351; // @[convert.scala 48:34]
  wire  _T_352; // @[convert.scala 49:36]
  wire [3:0] _T_354; // @[convert.scala 50:36]
  wire [3:0] _T_355; // @[convert.scala 50:36]
  wire [3:0] _T_356; // @[convert.scala 50:28]
  wire  _T_357; // @[convert.scala 51:31]
  wire  _T_358; // @[convert.scala 52:43]
  wire [9:0] _T_362; // @[Cat.scala 29:58]
  wire [3:0] _T_363; // @[Shift.scala 39:17]
  wire  _T_364; // @[Shift.scala 39:24]
  wire [1:0] _T_366; // @[Shift.scala 90:30]
  wire [7:0] _T_367; // @[Shift.scala 90:48]
  wire  _T_368; // @[Shift.scala 90:57]
  wire [1:0] _GEN_4; // @[Shift.scala 90:39]
  wire [1:0] _T_369; // @[Shift.scala 90:39]
  wire  _T_370; // @[Shift.scala 12:21]
  wire  _T_371; // @[Shift.scala 12:21]
  wire [7:0] _T_373; // @[Bitwise.scala 71:12]
  wire [9:0] _T_374; // @[Cat.scala 29:58]
  wire [9:0] _T_375; // @[Shift.scala 91:22]
  wire [2:0] _T_376; // @[Shift.scala 92:77]
  wire [5:0] _T_377; // @[Shift.scala 90:30]
  wire [3:0] _T_378; // @[Shift.scala 90:48]
  wire  _T_379; // @[Shift.scala 90:57]
  wire [5:0] _GEN_5; // @[Shift.scala 90:39]
  wire [5:0] _T_380; // @[Shift.scala 90:39]
  wire  _T_381; // @[Shift.scala 12:21]
  wire  _T_382; // @[Shift.scala 12:21]
  wire [3:0] _T_384; // @[Bitwise.scala 71:12]
  wire [9:0] _T_385; // @[Cat.scala 29:58]
  wire [9:0] _T_386; // @[Shift.scala 91:22]
  wire [1:0] _T_387; // @[Shift.scala 92:77]
  wire [7:0] _T_388; // @[Shift.scala 90:30]
  wire [1:0] _T_389; // @[Shift.scala 90:48]
  wire  _T_390; // @[Shift.scala 90:57]
  wire [7:0] _GEN_6; // @[Shift.scala 90:39]
  wire [7:0] _T_391; // @[Shift.scala 90:39]
  wire  _T_392; // @[Shift.scala 12:21]
  wire  _T_393; // @[Shift.scala 12:21]
  wire [1:0] _T_395; // @[Bitwise.scala 71:12]
  wire [9:0] _T_396; // @[Cat.scala 29:58]
  wire [9:0] _T_397; // @[Shift.scala 91:22]
  wire  _T_398; // @[Shift.scala 92:77]
  wire [8:0] _T_399; // @[Shift.scala 90:30]
  wire  _T_400; // @[Shift.scala 90:48]
  wire [8:0] _GEN_7; // @[Shift.scala 90:39]
  wire [8:0] _T_402; // @[Shift.scala 90:39]
  wire  _T_404; // @[Shift.scala 12:21]
  wire [9:0] _T_405; // @[Cat.scala 29:58]
  wire [9:0] _T_406; // @[Shift.scala 91:22]
  wire [9:0] _T_409; // @[Bitwise.scala 71:12]
  wire [9:0] _T_410; // @[Shift.scala 39:10]
  wire  _T_411; // @[convert.scala 55:31]
  wire  _T_412; // @[convert.scala 56:31]
  wire  _T_413; // @[convert.scala 57:31]
  wire  _T_414; // @[convert.scala 58:31]
  wire [6:0] _T_415; // @[convert.scala 59:69]
  wire  _T_416; // @[convert.scala 59:81]
  wire  _T_417; // @[convert.scala 59:50]
  wire  _T_419; // @[convert.scala 60:81]
  wire  _T_420; // @[convert.scala 61:44]
  wire  _T_421; // @[convert.scala 61:52]
  wire  _T_422; // @[convert.scala 61:36]
  wire  _T_423; // @[convert.scala 62:63]
  wire  _T_424; // @[convert.scala 62:103]
  wire  _T_425; // @[convert.scala 62:60]
  wire [6:0] _GEN_8; // @[convert.scala 63:56]
  wire [6:0] _T_428; // @[convert.scala 63:56]
  wire [7:0] _T_429; // @[Cat.scala 29:58]
  wire [7:0] _T_431; // @[Mux.scala 87:16]
  assign _T_1 = io_A[7]; // @[convert.scala 18:24]
  assign _T_2 = io_A[6]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[6:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[5:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[5:2]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[3:2]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8 != 2'h0; // @[LZD.scala 39:14]
  assign _T_10 = _T_8[1]; // @[LZD.scala 39:21]
  assign _T_11 = _T_8[0]; // @[LZD.scala 39:30]
  assign _T_12 = ~ _T_11; // @[LZD.scala 39:27]
  assign _T_13 = _T_10 | _T_12; // @[LZD.scala 39:25]
  assign _T_14 = {_T_9,_T_13}; // @[Cat.scala 29:58]
  assign _T_15 = _T_7[1:0]; // @[LZD.scala 44:32]
  assign _T_16 = _T_15 != 2'h0; // @[LZD.scala 39:14]
  assign _T_17 = _T_15[1]; // @[LZD.scala 39:21]
  assign _T_18 = _T_15[0]; // @[LZD.scala 39:30]
  assign _T_19 = ~ _T_18; // @[LZD.scala 39:27]
  assign _T_20 = _T_17 | _T_19; // @[LZD.scala 39:25]
  assign _T_21 = {_T_16,_T_20}; // @[Cat.scala 29:58]
  assign _T_22 = _T_14[1]; // @[Shift.scala 12:21]
  assign _T_23 = _T_21[1]; // @[Shift.scala 12:21]
  assign _T_24 = _T_22 | _T_23; // @[LZD.scala 49:16]
  assign _T_25 = ~ _T_23; // @[LZD.scala 49:27]
  assign _T_26 = _T_22 | _T_25; // @[LZD.scala 49:25]
  assign _T_27 = _T_14[0:0]; // @[LZD.scala 49:47]
  assign _T_28 = _T_21[0:0]; // @[LZD.scala 49:59]
  assign _T_29 = _T_22 ? _T_27 : _T_28; // @[LZD.scala 49:35]
  assign _T_31 = {_T_24,_T_26,_T_29}; // @[Cat.scala 29:58]
  assign _T_32 = _T_6[1:0]; // @[LZD.scala 44:32]
  assign _T_33 = _T_32 != 2'h0; // @[LZD.scala 39:14]
  assign _T_34 = _T_32[1]; // @[LZD.scala 39:21]
  assign _T_35 = _T_32[0]; // @[LZD.scala 39:30]
  assign _T_36 = ~ _T_35; // @[LZD.scala 39:27]
  assign _T_37 = _T_34 | _T_36; // @[LZD.scala 39:25]
  assign _T_38 = {_T_33,_T_37}; // @[Cat.scala 29:58]
  assign _T_39 = _T_31[2]; // @[Shift.scala 12:21]
  assign _T_41 = _T_31[1:0]; // @[LZD.scala 55:32]
  assign _T_42 = _T_39 ? _T_41 : _T_38; // @[LZD.scala 55:20]
  assign _T_43 = {_T_39,_T_42}; // @[Cat.scala 29:58]
  assign _T_44 = ~ _T_43; // @[convert.scala 21:22]
  assign _T_45 = io_A[4:0]; // @[convert.scala 22:36]
  assign _T_46 = _T_44 < 3'h5; // @[Shift.scala 16:24]
  assign _T_48 = _T_44[2]; // @[Shift.scala 12:21]
  assign _T_49 = _T_45[0:0]; // @[Shift.scala 64:52]
  assign _T_51 = {_T_49,4'h0}; // @[Cat.scala 29:58]
  assign _T_52 = _T_48 ? _T_51 : _T_45; // @[Shift.scala 64:27]
  assign _T_53 = _T_44[1:0]; // @[Shift.scala 66:70]
  assign _T_54 = _T_53[1]; // @[Shift.scala 12:21]
  assign _T_55 = _T_52[2:0]; // @[Shift.scala 64:52]
  assign _T_57 = {_T_55,2'h0}; // @[Cat.scala 29:58]
  assign _T_58 = _T_54 ? _T_57 : _T_52; // @[Shift.scala 64:27]
  assign _T_59 = _T_53[0:0]; // @[Shift.scala 66:70]
  assign _T_61 = _T_58[3:0]; // @[Shift.scala 64:52]
  assign _T_62 = {_T_61,1'h0}; // @[Cat.scala 29:58]
  assign _T_63 = _T_59 ? _T_62 : _T_58; // @[Shift.scala 64:27]
  assign _T_64 = _T_46 ? _T_63 : 5'h0; // @[Shift.scala 16:10]
  assign _T_65 = _T_64[4:4]; // @[convert.scala 23:34]
  assign decA_fraction = _T_64[3:0]; // @[convert.scala 24:34]
  assign _T_67 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_69 = _T_3 ? _T_44 : _T_43; // @[convert.scala 25:42]
  assign _T_72 = ~ _T_65; // @[convert.scala 26:67]
  assign _T_73 = _T_1 ? _T_72 : _T_65; // @[convert.scala 26:51]
  assign _T_74 = {_T_67,_T_69,_T_73}; // @[Cat.scala 29:58]
  assign _T_76 = io_A[6:0]; // @[convert.scala 29:56]
  assign _T_77 = _T_76 != 7'h0; // @[convert.scala 29:60]
  assign _T_78 = ~ _T_77; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_78; // @[convert.scala 29:39]
  assign _T_81 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_81 & _T_78; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_74); // @[convert.scala 32:24]
  assign _T_90 = io_B[7]; // @[convert.scala 18:24]
  assign _T_91 = io_B[6]; // @[convert.scala 18:40]
  assign _T_92 = _T_90 ^ _T_91; // @[convert.scala 18:36]
  assign _T_93 = io_B[6:1]; // @[convert.scala 19:24]
  assign _T_94 = io_B[5:0]; // @[convert.scala 19:43]
  assign _T_95 = _T_93 ^ _T_94; // @[convert.scala 19:39]
  assign _T_96 = _T_95[5:2]; // @[LZD.scala 43:32]
  assign _T_97 = _T_96[3:2]; // @[LZD.scala 43:32]
  assign _T_98 = _T_97 != 2'h0; // @[LZD.scala 39:14]
  assign _T_99 = _T_97[1]; // @[LZD.scala 39:21]
  assign _T_100 = _T_97[0]; // @[LZD.scala 39:30]
  assign _T_101 = ~ _T_100; // @[LZD.scala 39:27]
  assign _T_102 = _T_99 | _T_101; // @[LZD.scala 39:25]
  assign _T_103 = {_T_98,_T_102}; // @[Cat.scala 29:58]
  assign _T_104 = _T_96[1:0]; // @[LZD.scala 44:32]
  assign _T_105 = _T_104 != 2'h0; // @[LZD.scala 39:14]
  assign _T_106 = _T_104[1]; // @[LZD.scala 39:21]
  assign _T_107 = _T_104[0]; // @[LZD.scala 39:30]
  assign _T_108 = ~ _T_107; // @[LZD.scala 39:27]
  assign _T_109 = _T_106 | _T_108; // @[LZD.scala 39:25]
  assign _T_110 = {_T_105,_T_109}; // @[Cat.scala 29:58]
  assign _T_111 = _T_103[1]; // @[Shift.scala 12:21]
  assign _T_112 = _T_110[1]; // @[Shift.scala 12:21]
  assign _T_113 = _T_111 | _T_112; // @[LZD.scala 49:16]
  assign _T_114 = ~ _T_112; // @[LZD.scala 49:27]
  assign _T_115 = _T_111 | _T_114; // @[LZD.scala 49:25]
  assign _T_116 = _T_103[0:0]; // @[LZD.scala 49:47]
  assign _T_117 = _T_110[0:0]; // @[LZD.scala 49:59]
  assign _T_118 = _T_111 ? _T_116 : _T_117; // @[LZD.scala 49:35]
  assign _T_120 = {_T_113,_T_115,_T_118}; // @[Cat.scala 29:58]
  assign _T_121 = _T_95[1:0]; // @[LZD.scala 44:32]
  assign _T_122 = _T_121 != 2'h0; // @[LZD.scala 39:14]
  assign _T_123 = _T_121[1]; // @[LZD.scala 39:21]
  assign _T_124 = _T_121[0]; // @[LZD.scala 39:30]
  assign _T_125 = ~ _T_124; // @[LZD.scala 39:27]
  assign _T_126 = _T_123 | _T_125; // @[LZD.scala 39:25]
  assign _T_127 = {_T_122,_T_126}; // @[Cat.scala 29:58]
  assign _T_128 = _T_120[2]; // @[Shift.scala 12:21]
  assign _T_130 = _T_120[1:0]; // @[LZD.scala 55:32]
  assign _T_131 = _T_128 ? _T_130 : _T_127; // @[LZD.scala 55:20]
  assign _T_132 = {_T_128,_T_131}; // @[Cat.scala 29:58]
  assign _T_133 = ~ _T_132; // @[convert.scala 21:22]
  assign _T_134 = io_B[4:0]; // @[convert.scala 22:36]
  assign _T_135 = _T_133 < 3'h5; // @[Shift.scala 16:24]
  assign _T_137 = _T_133[2]; // @[Shift.scala 12:21]
  assign _T_138 = _T_134[0:0]; // @[Shift.scala 64:52]
  assign _T_140 = {_T_138,4'h0}; // @[Cat.scala 29:58]
  assign _T_141 = _T_137 ? _T_140 : _T_134; // @[Shift.scala 64:27]
  assign _T_142 = _T_133[1:0]; // @[Shift.scala 66:70]
  assign _T_143 = _T_142[1]; // @[Shift.scala 12:21]
  assign _T_144 = _T_141[2:0]; // @[Shift.scala 64:52]
  assign _T_146 = {_T_144,2'h0}; // @[Cat.scala 29:58]
  assign _T_147 = _T_143 ? _T_146 : _T_141; // @[Shift.scala 64:27]
  assign _T_148 = _T_142[0:0]; // @[Shift.scala 66:70]
  assign _T_150 = _T_147[3:0]; // @[Shift.scala 64:52]
  assign _T_151 = {_T_150,1'h0}; // @[Cat.scala 29:58]
  assign _T_152 = _T_148 ? _T_151 : _T_147; // @[Shift.scala 64:27]
  assign _T_153 = _T_135 ? _T_152 : 5'h0; // @[Shift.scala 16:10]
  assign _T_154 = _T_153[4:4]; // @[convert.scala 23:34]
  assign decB_fraction = _T_153[3:0]; // @[convert.scala 24:34]
  assign _T_156 = _T_92 == 1'h0; // @[convert.scala 25:26]
  assign _T_158 = _T_92 ? _T_133 : _T_132; // @[convert.scala 25:42]
  assign _T_161 = ~ _T_154; // @[convert.scala 26:67]
  assign _T_162 = _T_90 ? _T_161 : _T_154; // @[convert.scala 26:51]
  assign _T_163 = {_T_156,_T_158,_T_162}; // @[Cat.scala 29:58]
  assign _T_165 = io_B[6:0]; // @[convert.scala 29:56]
  assign _T_166 = _T_165 != 7'h0; // @[convert.scala 29:60]
  assign _T_167 = ~ _T_166; // @[convert.scala 29:41]
  assign decB_isNaR = _T_90 & _T_167; // @[convert.scala 29:39]
  assign _T_170 = _T_90 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_170 & _T_167; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_163); // @[convert.scala 32:24]
  assign aGTb = $signed(decA_scale) > $signed(decB_scale); // @[PositAdder.scala 24:32]
  assign greaterSign = aGTb ? _T_1 : _T_90; // @[PositAdder.scala 25:24]
  assign smallerSign = aGTb ? _T_90 : _T_1; // @[PositAdder.scala 26:24]
  assign greaterExp = aGTb ? $signed(decA_scale) : $signed(decB_scale); // @[PositAdder.scala 27:24]
  assign smallerExp = aGTb ? $signed(decB_scale) : $signed(decA_scale); // @[PositAdder.scala 28:24]
  assign greaterFrac = aGTb ? decA_fraction : decB_fraction; // @[PositAdder.scala 29:24]
  assign smallerFrac = aGTb ? decB_fraction : decA_fraction; // @[PositAdder.scala 30:24]
  assign smallerZero = aGTb ? decB_isZero : decA_isZero; // @[PositAdder.scala 31:24]
  assign _T_179 = $signed(greaterExp) - $signed(smallerExp); // @[PositAdder.scala 32:32]
  assign scale_diff = $signed(_T_179); // @[PositAdder.scala 32:32]
  assign _T_180 = ~ greaterSign; // @[PositAdder.scala 33:38]
  assign greaterSig = {greaterSign,_T_180,greaterFrac}; // @[Cat.scala 29:58]
  assign _T_182 = smallerSign | smallerZero; // @[PositAdder.scala 34:52]
  assign _T_183 = ~ _T_182; // @[PositAdder.scala 34:38]
  assign _T_186 = {smallerSign,_T_183,smallerFrac,3'h0}; // @[Cat.scala 29:58]
  assign _T_187 = $unsigned(scale_diff); // @[PositAdder.scala 35:68]
  assign _T_188 = _T_187 < 5'h9; // @[Shift.scala 39:24]
  assign _T_189 = _T_187[3:0]; // @[Shift.scala 40:44]
  assign _T_190 = _T_186[8:8]; // @[Shift.scala 90:30]
  assign _T_191 = _T_186[7:0]; // @[Shift.scala 90:48]
  assign _T_192 = _T_191 != 8'h0; // @[Shift.scala 90:57]
  assign _T_193 = _T_190 | _T_192; // @[Shift.scala 90:39]
  assign _T_194 = _T_189[3]; // @[Shift.scala 12:21]
  assign _T_195 = _T_186[8]; // @[Shift.scala 12:21]
  assign _T_197 = _T_195 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_198 = {_T_197,_T_193}; // @[Cat.scala 29:58]
  assign _T_199 = _T_194 ? _T_198 : _T_186; // @[Shift.scala 91:22]
  assign _T_200 = _T_189[2:0]; // @[Shift.scala 92:77]
  assign _T_201 = _T_199[8:4]; // @[Shift.scala 90:30]
  assign _T_202 = _T_199[3:0]; // @[Shift.scala 90:48]
  assign _T_203 = _T_202 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_0 = {{4'd0}, _T_203}; // @[Shift.scala 90:39]
  assign _T_204 = _T_201 | _GEN_0; // @[Shift.scala 90:39]
  assign _T_205 = _T_200[2]; // @[Shift.scala 12:21]
  assign _T_206 = _T_199[8]; // @[Shift.scala 12:21]
  assign _T_208 = _T_206 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_209 = {_T_208,_T_204}; // @[Cat.scala 29:58]
  assign _T_210 = _T_205 ? _T_209 : _T_199; // @[Shift.scala 91:22]
  assign _T_211 = _T_200[1:0]; // @[Shift.scala 92:77]
  assign _T_212 = _T_210[8:2]; // @[Shift.scala 90:30]
  assign _T_213 = _T_210[1:0]; // @[Shift.scala 90:48]
  assign _T_214 = _T_213 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_1 = {{6'd0}, _T_214}; // @[Shift.scala 90:39]
  assign _T_215 = _T_212 | _GEN_1; // @[Shift.scala 90:39]
  assign _T_216 = _T_211[1]; // @[Shift.scala 12:21]
  assign _T_217 = _T_210[8]; // @[Shift.scala 12:21]
  assign _T_219 = _T_217 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_220 = {_T_219,_T_215}; // @[Cat.scala 29:58]
  assign _T_221 = _T_216 ? _T_220 : _T_210; // @[Shift.scala 91:22]
  assign _T_222 = _T_211[0:0]; // @[Shift.scala 92:77]
  assign _T_223 = _T_221[8:1]; // @[Shift.scala 90:30]
  assign _T_224 = _T_221[0:0]; // @[Shift.scala 90:48]
  assign _GEN_2 = {{7'd0}, _T_224}; // @[Shift.scala 90:39]
  assign _T_226 = _T_223 | _GEN_2; // @[Shift.scala 90:39]
  assign _T_228 = _T_221[8]; // @[Shift.scala 12:21]
  assign _T_229 = {_T_228,_T_226}; // @[Cat.scala 29:58]
  assign _T_230 = _T_222 ? _T_229 : _T_221; // @[Shift.scala 91:22]
  assign _T_233 = _T_195 ? 9'h1ff : 9'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_188 ? _T_230 : _T_233; // @[Shift.scala 39:10]
  assign _T_234 = smallerSig[8:3]; // @[PositAdder.scala 36:45]
  assign rawSumSig = greaterSig + _T_234; // @[PositAdder.scala 36:32]
  assign _T_235 = _T_1 ^ _T_90; // @[PositAdder.scala 37:31]
  assign _T_236 = rawSumSig[6:6]; // @[PositAdder.scala 37:59]
  assign sumSign = _T_235 ^ _T_236; // @[PositAdder.scala 37:43]
  assign _T_237 = greaterSig + _T_234; // @[PositAdder.scala 38:48]
  assign _T_238 = smallerSig[2:0]; // @[PositAdder.scala 38:63]
  assign signSumSig = {sumSign,_T_237,_T_238}; // @[Cat.scala 29:58]
  assign _T_240 = signSumSig[9:1]; // @[PositAdder.scala 40:31]
  assign _T_241 = signSumSig[8:0]; // @[PositAdder.scala 40:66]
  assign sumXor = _T_240 ^ _T_241; // @[PositAdder.scala 40:49]
  assign _T_242 = sumXor[8:1]; // @[LZD.scala 43:32]
  assign _T_243 = _T_242[7:4]; // @[LZD.scala 43:32]
  assign _T_244 = _T_243[3:2]; // @[LZD.scala 43:32]
  assign _T_245 = _T_244 != 2'h0; // @[LZD.scala 39:14]
  assign _T_246 = _T_244[1]; // @[LZD.scala 39:21]
  assign _T_247 = _T_244[0]; // @[LZD.scala 39:30]
  assign _T_248 = ~ _T_247; // @[LZD.scala 39:27]
  assign _T_249 = _T_246 | _T_248; // @[LZD.scala 39:25]
  assign _T_250 = {_T_245,_T_249}; // @[Cat.scala 29:58]
  assign _T_251 = _T_243[1:0]; // @[LZD.scala 44:32]
  assign _T_252 = _T_251 != 2'h0; // @[LZD.scala 39:14]
  assign _T_253 = _T_251[1]; // @[LZD.scala 39:21]
  assign _T_254 = _T_251[0]; // @[LZD.scala 39:30]
  assign _T_255 = ~ _T_254; // @[LZD.scala 39:27]
  assign _T_256 = _T_253 | _T_255; // @[LZD.scala 39:25]
  assign _T_257 = {_T_252,_T_256}; // @[Cat.scala 29:58]
  assign _T_258 = _T_250[1]; // @[Shift.scala 12:21]
  assign _T_259 = _T_257[1]; // @[Shift.scala 12:21]
  assign _T_260 = _T_258 | _T_259; // @[LZD.scala 49:16]
  assign _T_261 = ~ _T_259; // @[LZD.scala 49:27]
  assign _T_262 = _T_258 | _T_261; // @[LZD.scala 49:25]
  assign _T_263 = _T_250[0:0]; // @[LZD.scala 49:47]
  assign _T_264 = _T_257[0:0]; // @[LZD.scala 49:59]
  assign _T_265 = _T_258 ? _T_263 : _T_264; // @[LZD.scala 49:35]
  assign _T_267 = {_T_260,_T_262,_T_265}; // @[Cat.scala 29:58]
  assign _T_268 = _T_242[3:0]; // @[LZD.scala 44:32]
  assign _T_269 = _T_268[3:2]; // @[LZD.scala 43:32]
  assign _T_270 = _T_269 != 2'h0; // @[LZD.scala 39:14]
  assign _T_271 = _T_269[1]; // @[LZD.scala 39:21]
  assign _T_272 = _T_269[0]; // @[LZD.scala 39:30]
  assign _T_273 = ~ _T_272; // @[LZD.scala 39:27]
  assign _T_274 = _T_271 | _T_273; // @[LZD.scala 39:25]
  assign _T_275 = {_T_270,_T_274}; // @[Cat.scala 29:58]
  assign _T_276 = _T_268[1:0]; // @[LZD.scala 44:32]
  assign _T_277 = _T_276 != 2'h0; // @[LZD.scala 39:14]
  assign _T_278 = _T_276[1]; // @[LZD.scala 39:21]
  assign _T_279 = _T_276[0]; // @[LZD.scala 39:30]
  assign _T_280 = ~ _T_279; // @[LZD.scala 39:27]
  assign _T_281 = _T_278 | _T_280; // @[LZD.scala 39:25]
  assign _T_282 = {_T_277,_T_281}; // @[Cat.scala 29:58]
  assign _T_283 = _T_275[1]; // @[Shift.scala 12:21]
  assign _T_284 = _T_282[1]; // @[Shift.scala 12:21]
  assign _T_285 = _T_283 | _T_284; // @[LZD.scala 49:16]
  assign _T_286 = ~ _T_284; // @[LZD.scala 49:27]
  assign _T_287 = _T_283 | _T_286; // @[LZD.scala 49:25]
  assign _T_288 = _T_275[0:0]; // @[LZD.scala 49:47]
  assign _T_289 = _T_282[0:0]; // @[LZD.scala 49:59]
  assign _T_290 = _T_283 ? _T_288 : _T_289; // @[LZD.scala 49:35]
  assign _T_292 = {_T_285,_T_287,_T_290}; // @[Cat.scala 29:58]
  assign _T_293 = _T_267[2]; // @[Shift.scala 12:21]
  assign _T_294 = _T_292[2]; // @[Shift.scala 12:21]
  assign _T_295 = _T_293 | _T_294; // @[LZD.scala 49:16]
  assign _T_296 = ~ _T_294; // @[LZD.scala 49:27]
  assign _T_297 = _T_293 | _T_296; // @[LZD.scala 49:25]
  assign _T_298 = _T_267[1:0]; // @[LZD.scala 49:47]
  assign _T_299 = _T_292[1:0]; // @[LZD.scala 49:59]
  assign _T_300 = _T_293 ? _T_298 : _T_299; // @[LZD.scala 49:35]
  assign _T_302 = {_T_295,_T_297,_T_300}; // @[Cat.scala 29:58]
  assign _T_303 = sumXor[0:0]; // @[LZD.scala 44:32]
  assign _T_305 = _T_302[3]; // @[Shift.scala 12:21]
  assign _T_308 = {2'h3,_T_303}; // @[Cat.scala 29:58]
  assign _T_309 = _T_302[2:0]; // @[LZD.scala 55:32]
  assign _T_310 = _T_305 ? _T_309 : _T_308; // @[LZD.scala 55:20]
  assign sumLZD = {_T_305,_T_310}; // @[Cat.scala 29:58]
  assign _T_311 = {1'h1,_T_305,_T_310}; // @[Cat.scala 29:58]
  assign _T_312 = $signed(_T_311); // @[PositAdder.scala 42:38]
  assign _T_314 = $signed(_T_312) + $signed(5'sh2); // @[PositAdder.scala 42:45]
  assign scaleBias = $signed(_T_314); // @[PositAdder.scala 42:45]
  assign sumScale = $signed(greaterExp) + $signed(scaleBias); // @[PositAdder.scala 43:32]
  assign overflow = $signed(sumScale) > $signed(6'shc); // @[PositAdder.scala 44:30]
  assign normalShift = ~ sumLZD; // @[PositAdder.scala 45:22]
  assign _T_315 = signSumSig[7:0]; // @[PositAdder.scala 46:36]
  assign _T_316 = normalShift < 4'h8; // @[Shift.scala 16:24]
  assign _T_317 = normalShift[2:0]; // @[Shift.scala 17:37]
  assign _T_318 = _T_317[2]; // @[Shift.scala 12:21]
  assign _T_319 = _T_315[3:0]; // @[Shift.scala 64:52]
  assign _T_321 = {_T_319,4'h0}; // @[Cat.scala 29:58]
  assign _T_322 = _T_318 ? _T_321 : _T_315; // @[Shift.scala 64:27]
  assign _T_323 = _T_317[1:0]; // @[Shift.scala 66:70]
  assign _T_324 = _T_323[1]; // @[Shift.scala 12:21]
  assign _T_325 = _T_322[5:0]; // @[Shift.scala 64:52]
  assign _T_327 = {_T_325,2'h0}; // @[Cat.scala 29:58]
  assign _T_328 = _T_324 ? _T_327 : _T_322; // @[Shift.scala 64:27]
  assign _T_329 = _T_323[0:0]; // @[Shift.scala 66:70]
  assign _T_331 = _T_328[6:0]; // @[Shift.scala 64:52]
  assign _T_332 = {_T_331,1'h0}; // @[Cat.scala 29:58]
  assign _T_333 = _T_329 ? _T_332 : _T_328; // @[Shift.scala 64:27]
  assign shiftSig = _T_316 ? _T_333 : 8'h0; // @[Shift.scala 16:10]
  assign _T_334 = overflow ? $signed(6'shc) : $signed(sumScale); // @[PositAdder.scala 51:24]
  assign decS_fraction = shiftSig[7:4]; // @[PositAdder.scala 52:34]
  assign decS_isNaR = decA_isNaR | decB_isNaR; // @[PositAdder.scala 53:32]
  assign _T_337 = signSumSig != 10'h0; // @[PositAdder.scala 54:33]
  assign _T_338 = ~ _T_337; // @[PositAdder.scala 54:21]
  assign _T_339 = decA_isZero & decB_isZero; // @[PositAdder.scala 54:52]
  assign decS_isZero = _T_338 | _T_339; // @[PositAdder.scala 54:37]
  assign _T_341 = shiftSig[3:2]; // @[PositAdder.scala 55:33]
  assign _T_342 = shiftSig[1]; // @[PositAdder.scala 55:49]
  assign _T_343 = shiftSig[0]; // @[PositAdder.scala 55:63]
  assign _T_344 = _T_342 | _T_343; // @[PositAdder.scala 55:53]
  assign _GEN_3 = _T_334[4:0]; // @[PositAdder.scala 48:25 PositAdder.scala 51:18]
  assign decS_scale = $signed(_GEN_3); // @[PositAdder.scala 48:25 PositAdder.scala 51:18]
  assign _T_347 = decS_scale[0]; // @[convert.scala 46:61]
  assign _T_348 = ~ _T_347; // @[convert.scala 46:52]
  assign _T_350 = sumSign ? _T_348 : _T_347; // @[convert.scala 46:42]
  assign _T_351 = decS_scale[4:1]; // @[convert.scala 48:34]
  assign _T_352 = _T_351[3:3]; // @[convert.scala 49:36]
  assign _T_354 = ~ _T_351; // @[convert.scala 50:36]
  assign _T_355 = $signed(_T_354); // @[convert.scala 50:36]
  assign _T_356 = _T_352 ? $signed(_T_355) : $signed(_T_351); // @[convert.scala 50:28]
  assign _T_357 = _T_352 ^ sumSign; // @[convert.scala 51:31]
  assign _T_358 = ~ _T_357; // @[convert.scala 52:43]
  assign _T_362 = {_T_358,_T_357,_T_350,decS_fraction,_T_341,_T_344}; // @[Cat.scala 29:58]
  assign _T_363 = $unsigned(_T_356); // @[Shift.scala 39:17]
  assign _T_364 = _T_363 < 4'ha; // @[Shift.scala 39:24]
  assign _T_366 = _T_362[9:8]; // @[Shift.scala 90:30]
  assign _T_367 = _T_362[7:0]; // @[Shift.scala 90:48]
  assign _T_368 = _T_367 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_4 = {{1'd0}, _T_368}; // @[Shift.scala 90:39]
  assign _T_369 = _T_366 | _GEN_4; // @[Shift.scala 90:39]
  assign _T_370 = _T_363[3]; // @[Shift.scala 12:21]
  assign _T_371 = _T_362[9]; // @[Shift.scala 12:21]
  assign _T_373 = _T_371 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_374 = {_T_373,_T_369}; // @[Cat.scala 29:58]
  assign _T_375 = _T_370 ? _T_374 : _T_362; // @[Shift.scala 91:22]
  assign _T_376 = _T_363[2:0]; // @[Shift.scala 92:77]
  assign _T_377 = _T_375[9:4]; // @[Shift.scala 90:30]
  assign _T_378 = _T_375[3:0]; // @[Shift.scala 90:48]
  assign _T_379 = _T_378 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_5 = {{5'd0}, _T_379}; // @[Shift.scala 90:39]
  assign _T_380 = _T_377 | _GEN_5; // @[Shift.scala 90:39]
  assign _T_381 = _T_376[2]; // @[Shift.scala 12:21]
  assign _T_382 = _T_375[9]; // @[Shift.scala 12:21]
  assign _T_384 = _T_382 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_385 = {_T_384,_T_380}; // @[Cat.scala 29:58]
  assign _T_386 = _T_381 ? _T_385 : _T_375; // @[Shift.scala 91:22]
  assign _T_387 = _T_376[1:0]; // @[Shift.scala 92:77]
  assign _T_388 = _T_386[9:2]; // @[Shift.scala 90:30]
  assign _T_389 = _T_386[1:0]; // @[Shift.scala 90:48]
  assign _T_390 = _T_389 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_6 = {{7'd0}, _T_390}; // @[Shift.scala 90:39]
  assign _T_391 = _T_388 | _GEN_6; // @[Shift.scala 90:39]
  assign _T_392 = _T_387[1]; // @[Shift.scala 12:21]
  assign _T_393 = _T_386[9]; // @[Shift.scala 12:21]
  assign _T_395 = _T_393 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_396 = {_T_395,_T_391}; // @[Cat.scala 29:58]
  assign _T_397 = _T_392 ? _T_396 : _T_386; // @[Shift.scala 91:22]
  assign _T_398 = _T_387[0:0]; // @[Shift.scala 92:77]
  assign _T_399 = _T_397[9:1]; // @[Shift.scala 90:30]
  assign _T_400 = _T_397[0:0]; // @[Shift.scala 90:48]
  assign _GEN_7 = {{8'd0}, _T_400}; // @[Shift.scala 90:39]
  assign _T_402 = _T_399 | _GEN_7; // @[Shift.scala 90:39]
  assign _T_404 = _T_397[9]; // @[Shift.scala 12:21]
  assign _T_405 = {_T_404,_T_402}; // @[Cat.scala 29:58]
  assign _T_406 = _T_398 ? _T_405 : _T_397; // @[Shift.scala 91:22]
  assign _T_409 = _T_371 ? 10'h3ff : 10'h0; // @[Bitwise.scala 71:12]
  assign _T_410 = _T_364 ? _T_406 : _T_409; // @[Shift.scala 39:10]
  assign _T_411 = _T_410[3]; // @[convert.scala 55:31]
  assign _T_412 = _T_410[2]; // @[convert.scala 56:31]
  assign _T_413 = _T_410[1]; // @[convert.scala 57:31]
  assign _T_414 = _T_410[0]; // @[convert.scala 58:31]
  assign _T_415 = _T_410[9:3]; // @[convert.scala 59:69]
  assign _T_416 = _T_415 != 7'h0; // @[convert.scala 59:81]
  assign _T_417 = ~ _T_416; // @[convert.scala 59:50]
  assign _T_419 = _T_415 == 7'h7f; // @[convert.scala 60:81]
  assign _T_420 = _T_411 | _T_413; // @[convert.scala 61:44]
  assign _T_421 = _T_420 | _T_414; // @[convert.scala 61:52]
  assign _T_422 = _T_412 & _T_421; // @[convert.scala 61:36]
  assign _T_423 = ~ _T_419; // @[convert.scala 62:63]
  assign _T_424 = _T_423 & _T_422; // @[convert.scala 62:103]
  assign _T_425 = _T_417 | _T_424; // @[convert.scala 62:60]
  assign _GEN_8 = {{6'd0}, _T_425}; // @[convert.scala 63:56]
  assign _T_428 = _T_415 + _GEN_8; // @[convert.scala 63:56]
  assign _T_429 = {sumSign,_T_428}; // @[Cat.scala 29:58]
  assign _T_431 = decS_isZero ? 8'h0 : _T_429; // @[Mux.scala 87:16]
  assign io_S = decS_isNaR ? 8'h80 : _T_431; // @[PositAdder.scala 57:8]
endmodule
