module PositAdder12_1(
  input         clock,
  input         reset,
  input  [11:0] io_A,
  input  [11:0] io_B,
  output [11:0] io_S
);
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [9:0] _T_4; // @[convert.scala 19:24]
  wire [9:0] _T_5; // @[convert.scala 19:43]
  wire [9:0] _T_6; // @[convert.scala 19:39]
  wire [7:0] _T_7; // @[LZD.scala 43:32]
  wire [3:0] _T_8; // @[LZD.scala 43:32]
  wire [1:0] _T_9; // @[LZD.scala 43:32]
  wire  _T_10; // @[LZD.scala 39:14]
  wire  _T_11; // @[LZD.scala 39:21]
  wire  _T_12; // @[LZD.scala 39:30]
  wire  _T_13; // @[LZD.scala 39:27]
  wire  _T_14; // @[LZD.scala 39:25]
  wire [1:0] _T_15; // @[Cat.scala 29:58]
  wire [1:0] _T_16; // @[LZD.scala 44:32]
  wire  _T_17; // @[LZD.scala 39:14]
  wire  _T_18; // @[LZD.scala 39:21]
  wire  _T_19; // @[LZD.scala 39:30]
  wire  _T_20; // @[LZD.scala 39:27]
  wire  _T_21; // @[LZD.scala 39:25]
  wire [1:0] _T_22; // @[Cat.scala 29:58]
  wire  _T_23; // @[Shift.scala 12:21]
  wire  _T_24; // @[Shift.scala 12:21]
  wire  _T_25; // @[LZD.scala 49:16]
  wire  _T_26; // @[LZD.scala 49:27]
  wire  _T_27; // @[LZD.scala 49:25]
  wire  _T_28; // @[LZD.scala 49:47]
  wire  _T_29; // @[LZD.scala 49:59]
  wire  _T_30; // @[LZD.scala 49:35]
  wire [2:0] _T_32; // @[Cat.scala 29:58]
  wire [3:0] _T_33; // @[LZD.scala 44:32]
  wire [1:0] _T_34; // @[LZD.scala 43:32]
  wire  _T_35; // @[LZD.scala 39:14]
  wire  _T_36; // @[LZD.scala 39:21]
  wire  _T_37; // @[LZD.scala 39:30]
  wire  _T_38; // @[LZD.scala 39:27]
  wire  _T_39; // @[LZD.scala 39:25]
  wire [1:0] _T_40; // @[Cat.scala 29:58]
  wire [1:0] _T_41; // @[LZD.scala 44:32]
  wire  _T_42; // @[LZD.scala 39:14]
  wire  _T_43; // @[LZD.scala 39:21]
  wire  _T_44; // @[LZD.scala 39:30]
  wire  _T_45; // @[LZD.scala 39:27]
  wire  _T_46; // @[LZD.scala 39:25]
  wire [1:0] _T_47; // @[Cat.scala 29:58]
  wire  _T_48; // @[Shift.scala 12:21]
  wire  _T_49; // @[Shift.scala 12:21]
  wire  _T_50; // @[LZD.scala 49:16]
  wire  _T_51; // @[LZD.scala 49:27]
  wire  _T_52; // @[LZD.scala 49:25]
  wire  _T_53; // @[LZD.scala 49:47]
  wire  _T_54; // @[LZD.scala 49:59]
  wire  _T_55; // @[LZD.scala 49:35]
  wire [2:0] _T_57; // @[Cat.scala 29:58]
  wire  _T_58; // @[Shift.scala 12:21]
  wire  _T_59; // @[Shift.scala 12:21]
  wire  _T_60; // @[LZD.scala 49:16]
  wire  _T_61; // @[LZD.scala 49:27]
  wire  _T_62; // @[LZD.scala 49:25]
  wire [1:0] _T_63; // @[LZD.scala 49:47]
  wire [1:0] _T_64; // @[LZD.scala 49:59]
  wire [1:0] _T_65; // @[LZD.scala 49:35]
  wire [3:0] _T_67; // @[Cat.scala 29:58]
  wire [1:0] _T_68; // @[LZD.scala 44:32]
  wire  _T_69; // @[LZD.scala 39:14]
  wire  _T_70; // @[LZD.scala 39:21]
  wire  _T_71; // @[LZD.scala 39:30]
  wire  _T_72; // @[LZD.scala 39:27]
  wire  _T_73; // @[LZD.scala 39:25]
  wire  _T_75; // @[Shift.scala 12:21]
  wire [2:0] _T_77; // @[Cat.scala 29:58]
  wire [2:0] _T_78; // @[LZD.scala 55:32]
  wire [2:0] _T_79; // @[LZD.scala 55:20]
  wire [3:0] _T_80; // @[Cat.scala 29:58]
  wire [3:0] _T_81; // @[convert.scala 21:22]
  wire [8:0] _T_82; // @[convert.scala 22:36]
  wire  _T_83; // @[Shift.scala 16:24]
  wire  _T_85; // @[Shift.scala 12:21]
  wire  _T_86; // @[Shift.scala 64:52]
  wire [8:0] _T_88; // @[Cat.scala 29:58]
  wire [8:0] _T_89; // @[Shift.scala 64:27]
  wire [2:0] _T_90; // @[Shift.scala 66:70]
  wire  _T_91; // @[Shift.scala 12:21]
  wire [4:0] _T_92; // @[Shift.scala 64:52]
  wire [8:0] _T_94; // @[Cat.scala 29:58]
  wire [8:0] _T_95; // @[Shift.scala 64:27]
  wire [1:0] _T_96; // @[Shift.scala 66:70]
  wire  _T_97; // @[Shift.scala 12:21]
  wire [6:0] _T_98; // @[Shift.scala 64:52]
  wire [8:0] _T_100; // @[Cat.scala 29:58]
  wire [8:0] _T_101; // @[Shift.scala 64:27]
  wire  _T_102; // @[Shift.scala 66:70]
  wire [7:0] _T_104; // @[Shift.scala 64:52]
  wire [8:0] _T_105; // @[Cat.scala 29:58]
  wire [8:0] _T_106; // @[Shift.scala 64:27]
  wire [8:0] _T_107; // @[Shift.scala 16:10]
  wire  _T_108; // @[convert.scala 23:34]
  wire [7:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_110; // @[convert.scala 25:26]
  wire [3:0] _T_112; // @[convert.scala 25:42]
  wire  _T_115; // @[convert.scala 26:67]
  wire  _T_116; // @[convert.scala 26:51]
  wire [5:0] _T_117; // @[Cat.scala 29:58]
  wire [10:0] _T_119; // @[convert.scala 29:56]
  wire  _T_120; // @[convert.scala 29:60]
  wire  _T_121; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_124; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [5:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_133; // @[convert.scala 18:24]
  wire  _T_134; // @[convert.scala 18:40]
  wire  _T_135; // @[convert.scala 18:36]
  wire [9:0] _T_136; // @[convert.scala 19:24]
  wire [9:0] _T_137; // @[convert.scala 19:43]
  wire [9:0] _T_138; // @[convert.scala 19:39]
  wire [7:0] _T_139; // @[LZD.scala 43:32]
  wire [3:0] _T_140; // @[LZD.scala 43:32]
  wire [1:0] _T_141; // @[LZD.scala 43:32]
  wire  _T_142; // @[LZD.scala 39:14]
  wire  _T_143; // @[LZD.scala 39:21]
  wire  _T_144; // @[LZD.scala 39:30]
  wire  _T_145; // @[LZD.scala 39:27]
  wire  _T_146; // @[LZD.scala 39:25]
  wire [1:0] _T_147; // @[Cat.scala 29:58]
  wire [1:0] _T_148; // @[LZD.scala 44:32]
  wire  _T_149; // @[LZD.scala 39:14]
  wire  _T_150; // @[LZD.scala 39:21]
  wire  _T_151; // @[LZD.scala 39:30]
  wire  _T_152; // @[LZD.scala 39:27]
  wire  _T_153; // @[LZD.scala 39:25]
  wire [1:0] _T_154; // @[Cat.scala 29:58]
  wire  _T_155; // @[Shift.scala 12:21]
  wire  _T_156; // @[Shift.scala 12:21]
  wire  _T_157; // @[LZD.scala 49:16]
  wire  _T_158; // @[LZD.scala 49:27]
  wire  _T_159; // @[LZD.scala 49:25]
  wire  _T_160; // @[LZD.scala 49:47]
  wire  _T_161; // @[LZD.scala 49:59]
  wire  _T_162; // @[LZD.scala 49:35]
  wire [2:0] _T_164; // @[Cat.scala 29:58]
  wire [3:0] _T_165; // @[LZD.scala 44:32]
  wire [1:0] _T_166; // @[LZD.scala 43:32]
  wire  _T_167; // @[LZD.scala 39:14]
  wire  _T_168; // @[LZD.scala 39:21]
  wire  _T_169; // @[LZD.scala 39:30]
  wire  _T_170; // @[LZD.scala 39:27]
  wire  _T_171; // @[LZD.scala 39:25]
  wire [1:0] _T_172; // @[Cat.scala 29:58]
  wire [1:0] _T_173; // @[LZD.scala 44:32]
  wire  _T_174; // @[LZD.scala 39:14]
  wire  _T_175; // @[LZD.scala 39:21]
  wire  _T_176; // @[LZD.scala 39:30]
  wire  _T_177; // @[LZD.scala 39:27]
  wire  _T_178; // @[LZD.scala 39:25]
  wire [1:0] _T_179; // @[Cat.scala 29:58]
  wire  _T_180; // @[Shift.scala 12:21]
  wire  _T_181; // @[Shift.scala 12:21]
  wire  _T_182; // @[LZD.scala 49:16]
  wire  _T_183; // @[LZD.scala 49:27]
  wire  _T_184; // @[LZD.scala 49:25]
  wire  _T_185; // @[LZD.scala 49:47]
  wire  _T_186; // @[LZD.scala 49:59]
  wire  _T_187; // @[LZD.scala 49:35]
  wire [2:0] _T_189; // @[Cat.scala 29:58]
  wire  _T_190; // @[Shift.scala 12:21]
  wire  _T_191; // @[Shift.scala 12:21]
  wire  _T_192; // @[LZD.scala 49:16]
  wire  _T_193; // @[LZD.scala 49:27]
  wire  _T_194; // @[LZD.scala 49:25]
  wire [1:0] _T_195; // @[LZD.scala 49:47]
  wire [1:0] _T_196; // @[LZD.scala 49:59]
  wire [1:0] _T_197; // @[LZD.scala 49:35]
  wire [3:0] _T_199; // @[Cat.scala 29:58]
  wire [1:0] _T_200; // @[LZD.scala 44:32]
  wire  _T_201; // @[LZD.scala 39:14]
  wire  _T_202; // @[LZD.scala 39:21]
  wire  _T_203; // @[LZD.scala 39:30]
  wire  _T_204; // @[LZD.scala 39:27]
  wire  _T_205; // @[LZD.scala 39:25]
  wire  _T_207; // @[Shift.scala 12:21]
  wire [2:0] _T_209; // @[Cat.scala 29:58]
  wire [2:0] _T_210; // @[LZD.scala 55:32]
  wire [2:0] _T_211; // @[LZD.scala 55:20]
  wire [3:0] _T_212; // @[Cat.scala 29:58]
  wire [3:0] _T_213; // @[convert.scala 21:22]
  wire [8:0] _T_214; // @[convert.scala 22:36]
  wire  _T_215; // @[Shift.scala 16:24]
  wire  _T_217; // @[Shift.scala 12:21]
  wire  _T_218; // @[Shift.scala 64:52]
  wire [8:0] _T_220; // @[Cat.scala 29:58]
  wire [8:0] _T_221; // @[Shift.scala 64:27]
  wire [2:0] _T_222; // @[Shift.scala 66:70]
  wire  _T_223; // @[Shift.scala 12:21]
  wire [4:0] _T_224; // @[Shift.scala 64:52]
  wire [8:0] _T_226; // @[Cat.scala 29:58]
  wire [8:0] _T_227; // @[Shift.scala 64:27]
  wire [1:0] _T_228; // @[Shift.scala 66:70]
  wire  _T_229; // @[Shift.scala 12:21]
  wire [6:0] _T_230; // @[Shift.scala 64:52]
  wire [8:0] _T_232; // @[Cat.scala 29:58]
  wire [8:0] _T_233; // @[Shift.scala 64:27]
  wire  _T_234; // @[Shift.scala 66:70]
  wire [7:0] _T_236; // @[Shift.scala 64:52]
  wire [8:0] _T_237; // @[Cat.scala 29:58]
  wire [8:0] _T_238; // @[Shift.scala 64:27]
  wire [8:0] _T_239; // @[Shift.scala 16:10]
  wire  _T_240; // @[convert.scala 23:34]
  wire [7:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_242; // @[convert.scala 25:26]
  wire [3:0] _T_244; // @[convert.scala 25:42]
  wire  _T_247; // @[convert.scala 26:67]
  wire  _T_248; // @[convert.scala 26:51]
  wire [5:0] _T_249; // @[Cat.scala 29:58]
  wire [10:0] _T_251; // @[convert.scala 29:56]
  wire  _T_252; // @[convert.scala 29:60]
  wire  _T_253; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_256; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [5:0] decB_scale; // @[convert.scala 32:24]
  wire  aGTb; // @[PositAdder.scala 24:32]
  wire  greaterSign; // @[PositAdder.scala 25:24]
  wire  smallerSign; // @[PositAdder.scala 26:24]
  wire [5:0] greaterExp; // @[PositAdder.scala 27:24]
  wire [5:0] smallerExp; // @[PositAdder.scala 28:24]
  wire [7:0] greaterFrac; // @[PositAdder.scala 29:24]
  wire [7:0] smallerFrac; // @[PositAdder.scala 30:24]
  wire  smallerZero; // @[PositAdder.scala 31:24]
  wire [5:0] _T_265; // @[PositAdder.scala 32:32]
  wire [5:0] scale_diff; // @[PositAdder.scala 32:32]
  wire  _T_266; // @[PositAdder.scala 33:38]
  wire [9:0] greaterSig; // @[Cat.scala 29:58]
  wire  _T_268; // @[PositAdder.scala 34:52]
  wire  _T_269; // @[PositAdder.scala 34:38]
  wire [12:0] _T_272; // @[Cat.scala 29:58]
  wire [5:0] _T_273; // @[PositAdder.scala 35:68]
  wire  _T_274; // @[Shift.scala 39:24]
  wire [3:0] _T_275; // @[Shift.scala 40:44]
  wire [4:0] _T_276; // @[Shift.scala 90:30]
  wire [7:0] _T_277; // @[Shift.scala 90:48]
  wire  _T_278; // @[Shift.scala 90:57]
  wire [4:0] _GEN_0; // @[Shift.scala 90:39]
  wire [4:0] _T_279; // @[Shift.scala 90:39]
  wire  _T_280; // @[Shift.scala 12:21]
  wire  _T_281; // @[Shift.scala 12:21]
  wire [7:0] _T_283; // @[Bitwise.scala 71:12]
  wire [12:0] _T_284; // @[Cat.scala 29:58]
  wire [12:0] _T_285; // @[Shift.scala 91:22]
  wire [2:0] _T_286; // @[Shift.scala 92:77]
  wire [8:0] _T_287; // @[Shift.scala 90:30]
  wire [3:0] _T_288; // @[Shift.scala 90:48]
  wire  _T_289; // @[Shift.scala 90:57]
  wire [8:0] _GEN_1; // @[Shift.scala 90:39]
  wire [8:0] _T_290; // @[Shift.scala 90:39]
  wire  _T_291; // @[Shift.scala 12:21]
  wire  _T_292; // @[Shift.scala 12:21]
  wire [3:0] _T_294; // @[Bitwise.scala 71:12]
  wire [12:0] _T_295; // @[Cat.scala 29:58]
  wire [12:0] _T_296; // @[Shift.scala 91:22]
  wire [1:0] _T_297; // @[Shift.scala 92:77]
  wire [10:0] _T_298; // @[Shift.scala 90:30]
  wire [1:0] _T_299; // @[Shift.scala 90:48]
  wire  _T_300; // @[Shift.scala 90:57]
  wire [10:0] _GEN_2; // @[Shift.scala 90:39]
  wire [10:0] _T_301; // @[Shift.scala 90:39]
  wire  _T_302; // @[Shift.scala 12:21]
  wire  _T_303; // @[Shift.scala 12:21]
  wire [1:0] _T_305; // @[Bitwise.scala 71:12]
  wire [12:0] _T_306; // @[Cat.scala 29:58]
  wire [12:0] _T_307; // @[Shift.scala 91:22]
  wire  _T_308; // @[Shift.scala 92:77]
  wire [11:0] _T_309; // @[Shift.scala 90:30]
  wire  _T_310; // @[Shift.scala 90:48]
  wire [11:0] _GEN_3; // @[Shift.scala 90:39]
  wire [11:0] _T_312; // @[Shift.scala 90:39]
  wire  _T_314; // @[Shift.scala 12:21]
  wire [12:0] _T_315; // @[Cat.scala 29:58]
  wire [12:0] _T_316; // @[Shift.scala 91:22]
  wire [12:0] _T_319; // @[Bitwise.scala 71:12]
  wire [12:0] smallerSig; // @[Shift.scala 39:10]
  wire [9:0] _T_320; // @[PositAdder.scala 36:45]
  wire [10:0] rawSumSig; // @[PositAdder.scala 36:32]
  wire  _T_321; // @[PositAdder.scala 37:31]
  wire  _T_322; // @[PositAdder.scala 37:59]
  wire  sumSign; // @[PositAdder.scala 37:43]
  wire [9:0] _T_323; // @[PositAdder.scala 38:48]
  wire [2:0] _T_324; // @[PositAdder.scala 38:63]
  wire [13:0] signSumSig; // @[Cat.scala 29:58]
  wire [12:0] _T_326; // @[PositAdder.scala 40:31]
  wire [12:0] _T_327; // @[PositAdder.scala 40:66]
  wire [12:0] sumXor; // @[PositAdder.scala 40:49]
  wire [7:0] _T_328; // @[LZD.scala 43:32]
  wire [3:0] _T_329; // @[LZD.scala 43:32]
  wire [1:0] _T_330; // @[LZD.scala 43:32]
  wire  _T_331; // @[LZD.scala 39:14]
  wire  _T_332; // @[LZD.scala 39:21]
  wire  _T_333; // @[LZD.scala 39:30]
  wire  _T_334; // @[LZD.scala 39:27]
  wire  _T_335; // @[LZD.scala 39:25]
  wire [1:0] _T_336; // @[Cat.scala 29:58]
  wire [1:0] _T_337; // @[LZD.scala 44:32]
  wire  _T_338; // @[LZD.scala 39:14]
  wire  _T_339; // @[LZD.scala 39:21]
  wire  _T_340; // @[LZD.scala 39:30]
  wire  _T_341; // @[LZD.scala 39:27]
  wire  _T_342; // @[LZD.scala 39:25]
  wire [1:0] _T_343; // @[Cat.scala 29:58]
  wire  _T_344; // @[Shift.scala 12:21]
  wire  _T_345; // @[Shift.scala 12:21]
  wire  _T_346; // @[LZD.scala 49:16]
  wire  _T_347; // @[LZD.scala 49:27]
  wire  _T_348; // @[LZD.scala 49:25]
  wire  _T_349; // @[LZD.scala 49:47]
  wire  _T_350; // @[LZD.scala 49:59]
  wire  _T_351; // @[LZD.scala 49:35]
  wire [2:0] _T_353; // @[Cat.scala 29:58]
  wire [3:0] _T_354; // @[LZD.scala 44:32]
  wire [1:0] _T_355; // @[LZD.scala 43:32]
  wire  _T_356; // @[LZD.scala 39:14]
  wire  _T_357; // @[LZD.scala 39:21]
  wire  _T_358; // @[LZD.scala 39:30]
  wire  _T_359; // @[LZD.scala 39:27]
  wire  _T_360; // @[LZD.scala 39:25]
  wire [1:0] _T_361; // @[Cat.scala 29:58]
  wire [1:0] _T_362; // @[LZD.scala 44:32]
  wire  _T_363; // @[LZD.scala 39:14]
  wire  _T_364; // @[LZD.scala 39:21]
  wire  _T_365; // @[LZD.scala 39:30]
  wire  _T_366; // @[LZD.scala 39:27]
  wire  _T_367; // @[LZD.scala 39:25]
  wire [1:0] _T_368; // @[Cat.scala 29:58]
  wire  _T_369; // @[Shift.scala 12:21]
  wire  _T_370; // @[Shift.scala 12:21]
  wire  _T_371; // @[LZD.scala 49:16]
  wire  _T_372; // @[LZD.scala 49:27]
  wire  _T_373; // @[LZD.scala 49:25]
  wire  _T_374; // @[LZD.scala 49:47]
  wire  _T_375; // @[LZD.scala 49:59]
  wire  _T_376; // @[LZD.scala 49:35]
  wire [2:0] _T_378; // @[Cat.scala 29:58]
  wire  _T_379; // @[Shift.scala 12:21]
  wire  _T_380; // @[Shift.scala 12:21]
  wire  _T_381; // @[LZD.scala 49:16]
  wire  _T_382; // @[LZD.scala 49:27]
  wire  _T_383; // @[LZD.scala 49:25]
  wire [1:0] _T_384; // @[LZD.scala 49:47]
  wire [1:0] _T_385; // @[LZD.scala 49:59]
  wire [1:0] _T_386; // @[LZD.scala 49:35]
  wire [3:0] _T_388; // @[Cat.scala 29:58]
  wire [4:0] _T_389; // @[LZD.scala 44:32]
  wire [3:0] _T_390; // @[LZD.scala 43:32]
  wire [1:0] _T_391; // @[LZD.scala 43:32]
  wire  _T_392; // @[LZD.scala 39:14]
  wire  _T_393; // @[LZD.scala 39:21]
  wire  _T_394; // @[LZD.scala 39:30]
  wire  _T_395; // @[LZD.scala 39:27]
  wire  _T_396; // @[LZD.scala 39:25]
  wire [1:0] _T_397; // @[Cat.scala 29:58]
  wire [1:0] _T_398; // @[LZD.scala 44:32]
  wire  _T_399; // @[LZD.scala 39:14]
  wire  _T_400; // @[LZD.scala 39:21]
  wire  _T_401; // @[LZD.scala 39:30]
  wire  _T_402; // @[LZD.scala 39:27]
  wire  _T_403; // @[LZD.scala 39:25]
  wire [1:0] _T_404; // @[Cat.scala 29:58]
  wire  _T_405; // @[Shift.scala 12:21]
  wire  _T_406; // @[Shift.scala 12:21]
  wire  _T_407; // @[LZD.scala 49:16]
  wire  _T_408; // @[LZD.scala 49:27]
  wire  _T_409; // @[LZD.scala 49:25]
  wire  _T_410; // @[LZD.scala 49:47]
  wire  _T_411; // @[LZD.scala 49:59]
  wire  _T_412; // @[LZD.scala 49:35]
  wire [2:0] _T_414; // @[Cat.scala 29:58]
  wire  _T_415; // @[LZD.scala 44:32]
  wire  _T_417; // @[Shift.scala 12:21]
  wire [1:0] _T_419; // @[Cat.scala 29:58]
  wire [1:0] _T_420; // @[LZD.scala 55:32]
  wire [1:0] _T_421; // @[LZD.scala 55:20]
  wire [2:0] _T_422; // @[Cat.scala 29:58]
  wire  _T_423; // @[Shift.scala 12:21]
  wire [2:0] _T_425; // @[LZD.scala 55:32]
  wire [2:0] _T_426; // @[LZD.scala 55:20]
  wire [3:0] sumLZD; // @[Cat.scala 29:58]
  wire [4:0] _T_427; // @[Cat.scala 29:58]
  wire [4:0] _T_428; // @[PositAdder.scala 42:38]
  wire [4:0] _T_430; // @[PositAdder.scala 42:45]
  wire [4:0] scaleBias; // @[PositAdder.scala 42:45]
  wire [5:0] _GEN_4; // @[PositAdder.scala 43:32]
  wire [6:0] sumScale; // @[PositAdder.scala 43:32]
  wire  overflow; // @[PositAdder.scala 44:30]
  wire [3:0] normalShift; // @[PositAdder.scala 45:22]
  wire [11:0] _T_431; // @[PositAdder.scala 46:36]
  wire  _T_432; // @[Shift.scala 16:24]
  wire  _T_434; // @[Shift.scala 12:21]
  wire [3:0] _T_435; // @[Shift.scala 64:52]
  wire [11:0] _T_437; // @[Cat.scala 29:58]
  wire [11:0] _T_438; // @[Shift.scala 64:27]
  wire [2:0] _T_439; // @[Shift.scala 66:70]
  wire  _T_440; // @[Shift.scala 12:21]
  wire [7:0] _T_441; // @[Shift.scala 64:52]
  wire [11:0] _T_443; // @[Cat.scala 29:58]
  wire [11:0] _T_444; // @[Shift.scala 64:27]
  wire [1:0] _T_445; // @[Shift.scala 66:70]
  wire  _T_446; // @[Shift.scala 12:21]
  wire [9:0] _T_447; // @[Shift.scala 64:52]
  wire [11:0] _T_449; // @[Cat.scala 29:58]
  wire [11:0] _T_450; // @[Shift.scala 64:27]
  wire  _T_451; // @[Shift.scala 66:70]
  wire [10:0] _T_453; // @[Shift.scala 64:52]
  wire [11:0] _T_454; // @[Cat.scala 29:58]
  wire [11:0] _T_455; // @[Shift.scala 64:27]
  wire [11:0] shiftSig; // @[Shift.scala 16:10]
  wire [6:0] _T_456; // @[PositAdder.scala 51:24]
  wire [7:0] decS_fraction; // @[PositAdder.scala 52:34]
  wire  decS_isNaR; // @[PositAdder.scala 53:32]
  wire  _T_459; // @[PositAdder.scala 54:33]
  wire  _T_460; // @[PositAdder.scala 54:21]
  wire  _T_461; // @[PositAdder.scala 54:52]
  wire  decS_isZero; // @[PositAdder.scala 54:37]
  wire [1:0] _T_463; // @[PositAdder.scala 55:33]
  wire  _T_464; // @[PositAdder.scala 55:49]
  wire  _T_465; // @[PositAdder.scala 55:63]
  wire  _T_466; // @[PositAdder.scala 55:53]
  wire [5:0] _GEN_5; // @[PositAdder.scala 48:25 PositAdder.scala 51:18]
  wire [5:0] decS_scale; // @[PositAdder.scala 48:25 PositAdder.scala 51:18]
  wire  _T_469; // @[convert.scala 46:61]
  wire  _T_470; // @[convert.scala 46:52]
  wire  _T_472; // @[convert.scala 46:42]
  wire [4:0] _T_473; // @[convert.scala 48:34]
  wire  _T_474; // @[convert.scala 49:36]
  wire [4:0] _T_476; // @[convert.scala 50:36]
  wire [4:0] _T_477; // @[convert.scala 50:36]
  wire [4:0] _T_478; // @[convert.scala 50:28]
  wire  _T_479; // @[convert.scala 51:31]
  wire  _T_480; // @[convert.scala 52:43]
  wire [13:0] _T_484; // @[Cat.scala 29:58]
  wire [4:0] _T_485; // @[Shift.scala 39:17]
  wire  _T_486; // @[Shift.scala 39:24]
  wire [3:0] _T_487; // @[Shift.scala 40:44]
  wire [5:0] _T_488; // @[Shift.scala 90:30]
  wire [7:0] _T_489; // @[Shift.scala 90:48]
  wire  _T_490; // @[Shift.scala 90:57]
  wire [5:0] _GEN_6; // @[Shift.scala 90:39]
  wire [5:0] _T_491; // @[Shift.scala 90:39]
  wire  _T_492; // @[Shift.scala 12:21]
  wire  _T_493; // @[Shift.scala 12:21]
  wire [7:0] _T_495; // @[Bitwise.scala 71:12]
  wire [13:0] _T_496; // @[Cat.scala 29:58]
  wire [13:0] _T_497; // @[Shift.scala 91:22]
  wire [2:0] _T_498; // @[Shift.scala 92:77]
  wire [9:0] _T_499; // @[Shift.scala 90:30]
  wire [3:0] _T_500; // @[Shift.scala 90:48]
  wire  _T_501; // @[Shift.scala 90:57]
  wire [9:0] _GEN_7; // @[Shift.scala 90:39]
  wire [9:0] _T_502; // @[Shift.scala 90:39]
  wire  _T_503; // @[Shift.scala 12:21]
  wire  _T_504; // @[Shift.scala 12:21]
  wire [3:0] _T_506; // @[Bitwise.scala 71:12]
  wire [13:0] _T_507; // @[Cat.scala 29:58]
  wire [13:0] _T_508; // @[Shift.scala 91:22]
  wire [1:0] _T_509; // @[Shift.scala 92:77]
  wire [11:0] _T_510; // @[Shift.scala 90:30]
  wire [1:0] _T_511; // @[Shift.scala 90:48]
  wire  _T_512; // @[Shift.scala 90:57]
  wire [11:0] _GEN_8; // @[Shift.scala 90:39]
  wire [11:0] _T_513; // @[Shift.scala 90:39]
  wire  _T_514; // @[Shift.scala 12:21]
  wire  _T_515; // @[Shift.scala 12:21]
  wire [1:0] _T_517; // @[Bitwise.scala 71:12]
  wire [13:0] _T_518; // @[Cat.scala 29:58]
  wire [13:0] _T_519; // @[Shift.scala 91:22]
  wire  _T_520; // @[Shift.scala 92:77]
  wire [12:0] _T_521; // @[Shift.scala 90:30]
  wire  _T_522; // @[Shift.scala 90:48]
  wire [12:0] _GEN_9; // @[Shift.scala 90:39]
  wire [12:0] _T_524; // @[Shift.scala 90:39]
  wire  _T_526; // @[Shift.scala 12:21]
  wire [13:0] _T_527; // @[Cat.scala 29:58]
  wire [13:0] _T_528; // @[Shift.scala 91:22]
  wire [13:0] _T_531; // @[Bitwise.scala 71:12]
  wire [13:0] _T_532; // @[Shift.scala 39:10]
  wire  _T_533; // @[convert.scala 55:31]
  wire  _T_534; // @[convert.scala 56:31]
  wire  _T_535; // @[convert.scala 57:31]
  wire  _T_536; // @[convert.scala 58:31]
  wire [10:0] _T_537; // @[convert.scala 59:69]
  wire  _T_538; // @[convert.scala 59:81]
  wire  _T_539; // @[convert.scala 59:50]
  wire  _T_541; // @[convert.scala 60:81]
  wire  _T_542; // @[convert.scala 61:44]
  wire  _T_543; // @[convert.scala 61:52]
  wire  _T_544; // @[convert.scala 61:36]
  wire  _T_545; // @[convert.scala 62:63]
  wire  _T_546; // @[convert.scala 62:103]
  wire  _T_547; // @[convert.scala 62:60]
  wire [10:0] _GEN_10; // @[convert.scala 63:56]
  wire [10:0] _T_550; // @[convert.scala 63:56]
  wire [11:0] _T_551; // @[Cat.scala 29:58]
  wire [11:0] _T_553; // @[Mux.scala 87:16]
  assign _T_1 = io_A[11]; // @[convert.scala 18:24]
  assign _T_2 = io_A[10]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[10:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[9:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[9:2]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[7:4]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8[3:2]; // @[LZD.scala 43:32]
  assign _T_10 = _T_9 != 2'h0; // @[LZD.scala 39:14]
  assign _T_11 = _T_9[1]; // @[LZD.scala 39:21]
  assign _T_12 = _T_9[0]; // @[LZD.scala 39:30]
  assign _T_13 = ~ _T_12; // @[LZD.scala 39:27]
  assign _T_14 = _T_11 | _T_13; // @[LZD.scala 39:25]
  assign _T_15 = {_T_10,_T_14}; // @[Cat.scala 29:58]
  assign _T_16 = _T_8[1:0]; // @[LZD.scala 44:32]
  assign _T_17 = _T_16 != 2'h0; // @[LZD.scala 39:14]
  assign _T_18 = _T_16[1]; // @[LZD.scala 39:21]
  assign _T_19 = _T_16[0]; // @[LZD.scala 39:30]
  assign _T_20 = ~ _T_19; // @[LZD.scala 39:27]
  assign _T_21 = _T_18 | _T_20; // @[LZD.scala 39:25]
  assign _T_22 = {_T_17,_T_21}; // @[Cat.scala 29:58]
  assign _T_23 = _T_15[1]; // @[Shift.scala 12:21]
  assign _T_24 = _T_22[1]; // @[Shift.scala 12:21]
  assign _T_25 = _T_23 | _T_24; // @[LZD.scala 49:16]
  assign _T_26 = ~ _T_24; // @[LZD.scala 49:27]
  assign _T_27 = _T_23 | _T_26; // @[LZD.scala 49:25]
  assign _T_28 = _T_15[0:0]; // @[LZD.scala 49:47]
  assign _T_29 = _T_22[0:0]; // @[LZD.scala 49:59]
  assign _T_30 = _T_23 ? _T_28 : _T_29; // @[LZD.scala 49:35]
  assign _T_32 = {_T_25,_T_27,_T_30}; // @[Cat.scala 29:58]
  assign _T_33 = _T_7[3:0]; // @[LZD.scala 44:32]
  assign _T_34 = _T_33[3:2]; // @[LZD.scala 43:32]
  assign _T_35 = _T_34 != 2'h0; // @[LZD.scala 39:14]
  assign _T_36 = _T_34[1]; // @[LZD.scala 39:21]
  assign _T_37 = _T_34[0]; // @[LZD.scala 39:30]
  assign _T_38 = ~ _T_37; // @[LZD.scala 39:27]
  assign _T_39 = _T_36 | _T_38; // @[LZD.scala 39:25]
  assign _T_40 = {_T_35,_T_39}; // @[Cat.scala 29:58]
  assign _T_41 = _T_33[1:0]; // @[LZD.scala 44:32]
  assign _T_42 = _T_41 != 2'h0; // @[LZD.scala 39:14]
  assign _T_43 = _T_41[1]; // @[LZD.scala 39:21]
  assign _T_44 = _T_41[0]; // @[LZD.scala 39:30]
  assign _T_45 = ~ _T_44; // @[LZD.scala 39:27]
  assign _T_46 = _T_43 | _T_45; // @[LZD.scala 39:25]
  assign _T_47 = {_T_42,_T_46}; // @[Cat.scala 29:58]
  assign _T_48 = _T_40[1]; // @[Shift.scala 12:21]
  assign _T_49 = _T_47[1]; // @[Shift.scala 12:21]
  assign _T_50 = _T_48 | _T_49; // @[LZD.scala 49:16]
  assign _T_51 = ~ _T_49; // @[LZD.scala 49:27]
  assign _T_52 = _T_48 | _T_51; // @[LZD.scala 49:25]
  assign _T_53 = _T_40[0:0]; // @[LZD.scala 49:47]
  assign _T_54 = _T_47[0:0]; // @[LZD.scala 49:59]
  assign _T_55 = _T_48 ? _T_53 : _T_54; // @[LZD.scala 49:35]
  assign _T_57 = {_T_50,_T_52,_T_55}; // @[Cat.scala 29:58]
  assign _T_58 = _T_32[2]; // @[Shift.scala 12:21]
  assign _T_59 = _T_57[2]; // @[Shift.scala 12:21]
  assign _T_60 = _T_58 | _T_59; // @[LZD.scala 49:16]
  assign _T_61 = ~ _T_59; // @[LZD.scala 49:27]
  assign _T_62 = _T_58 | _T_61; // @[LZD.scala 49:25]
  assign _T_63 = _T_32[1:0]; // @[LZD.scala 49:47]
  assign _T_64 = _T_57[1:0]; // @[LZD.scala 49:59]
  assign _T_65 = _T_58 ? _T_63 : _T_64; // @[LZD.scala 49:35]
  assign _T_67 = {_T_60,_T_62,_T_65}; // @[Cat.scala 29:58]
  assign _T_68 = _T_6[1:0]; // @[LZD.scala 44:32]
  assign _T_69 = _T_68 != 2'h0; // @[LZD.scala 39:14]
  assign _T_70 = _T_68[1]; // @[LZD.scala 39:21]
  assign _T_71 = _T_68[0]; // @[LZD.scala 39:30]
  assign _T_72 = ~ _T_71; // @[LZD.scala 39:27]
  assign _T_73 = _T_70 | _T_72; // @[LZD.scala 39:25]
  assign _T_75 = _T_67[3]; // @[Shift.scala 12:21]
  assign _T_77 = {1'h1,_T_69,_T_73}; // @[Cat.scala 29:58]
  assign _T_78 = _T_67[2:0]; // @[LZD.scala 55:32]
  assign _T_79 = _T_75 ? _T_78 : _T_77; // @[LZD.scala 55:20]
  assign _T_80 = {_T_75,_T_79}; // @[Cat.scala 29:58]
  assign _T_81 = ~ _T_80; // @[convert.scala 21:22]
  assign _T_82 = io_A[8:0]; // @[convert.scala 22:36]
  assign _T_83 = _T_81 < 4'h9; // @[Shift.scala 16:24]
  assign _T_85 = _T_81[3]; // @[Shift.scala 12:21]
  assign _T_86 = _T_82[0:0]; // @[Shift.scala 64:52]
  assign _T_88 = {_T_86,8'h0}; // @[Cat.scala 29:58]
  assign _T_89 = _T_85 ? _T_88 : _T_82; // @[Shift.scala 64:27]
  assign _T_90 = _T_81[2:0]; // @[Shift.scala 66:70]
  assign _T_91 = _T_90[2]; // @[Shift.scala 12:21]
  assign _T_92 = _T_89[4:0]; // @[Shift.scala 64:52]
  assign _T_94 = {_T_92,4'h0}; // @[Cat.scala 29:58]
  assign _T_95 = _T_91 ? _T_94 : _T_89; // @[Shift.scala 64:27]
  assign _T_96 = _T_90[1:0]; // @[Shift.scala 66:70]
  assign _T_97 = _T_96[1]; // @[Shift.scala 12:21]
  assign _T_98 = _T_95[6:0]; // @[Shift.scala 64:52]
  assign _T_100 = {_T_98,2'h0}; // @[Cat.scala 29:58]
  assign _T_101 = _T_97 ? _T_100 : _T_95; // @[Shift.scala 64:27]
  assign _T_102 = _T_96[0:0]; // @[Shift.scala 66:70]
  assign _T_104 = _T_101[7:0]; // @[Shift.scala 64:52]
  assign _T_105 = {_T_104,1'h0}; // @[Cat.scala 29:58]
  assign _T_106 = _T_102 ? _T_105 : _T_101; // @[Shift.scala 64:27]
  assign _T_107 = _T_83 ? _T_106 : 9'h0; // @[Shift.scala 16:10]
  assign _T_108 = _T_107[8:8]; // @[convert.scala 23:34]
  assign decA_fraction = _T_107[7:0]; // @[convert.scala 24:34]
  assign _T_110 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_112 = _T_3 ? _T_81 : _T_80; // @[convert.scala 25:42]
  assign _T_115 = ~ _T_108; // @[convert.scala 26:67]
  assign _T_116 = _T_1 ? _T_115 : _T_108; // @[convert.scala 26:51]
  assign _T_117 = {_T_110,_T_112,_T_116}; // @[Cat.scala 29:58]
  assign _T_119 = io_A[10:0]; // @[convert.scala 29:56]
  assign _T_120 = _T_119 != 11'h0; // @[convert.scala 29:60]
  assign _T_121 = ~ _T_120; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_121; // @[convert.scala 29:39]
  assign _T_124 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_124 & _T_121; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_117); // @[convert.scala 32:24]
  assign _T_133 = io_B[11]; // @[convert.scala 18:24]
  assign _T_134 = io_B[10]; // @[convert.scala 18:40]
  assign _T_135 = _T_133 ^ _T_134; // @[convert.scala 18:36]
  assign _T_136 = io_B[10:1]; // @[convert.scala 19:24]
  assign _T_137 = io_B[9:0]; // @[convert.scala 19:43]
  assign _T_138 = _T_136 ^ _T_137; // @[convert.scala 19:39]
  assign _T_139 = _T_138[9:2]; // @[LZD.scala 43:32]
  assign _T_140 = _T_139[7:4]; // @[LZD.scala 43:32]
  assign _T_141 = _T_140[3:2]; // @[LZD.scala 43:32]
  assign _T_142 = _T_141 != 2'h0; // @[LZD.scala 39:14]
  assign _T_143 = _T_141[1]; // @[LZD.scala 39:21]
  assign _T_144 = _T_141[0]; // @[LZD.scala 39:30]
  assign _T_145 = ~ _T_144; // @[LZD.scala 39:27]
  assign _T_146 = _T_143 | _T_145; // @[LZD.scala 39:25]
  assign _T_147 = {_T_142,_T_146}; // @[Cat.scala 29:58]
  assign _T_148 = _T_140[1:0]; // @[LZD.scala 44:32]
  assign _T_149 = _T_148 != 2'h0; // @[LZD.scala 39:14]
  assign _T_150 = _T_148[1]; // @[LZD.scala 39:21]
  assign _T_151 = _T_148[0]; // @[LZD.scala 39:30]
  assign _T_152 = ~ _T_151; // @[LZD.scala 39:27]
  assign _T_153 = _T_150 | _T_152; // @[LZD.scala 39:25]
  assign _T_154 = {_T_149,_T_153}; // @[Cat.scala 29:58]
  assign _T_155 = _T_147[1]; // @[Shift.scala 12:21]
  assign _T_156 = _T_154[1]; // @[Shift.scala 12:21]
  assign _T_157 = _T_155 | _T_156; // @[LZD.scala 49:16]
  assign _T_158 = ~ _T_156; // @[LZD.scala 49:27]
  assign _T_159 = _T_155 | _T_158; // @[LZD.scala 49:25]
  assign _T_160 = _T_147[0:0]; // @[LZD.scala 49:47]
  assign _T_161 = _T_154[0:0]; // @[LZD.scala 49:59]
  assign _T_162 = _T_155 ? _T_160 : _T_161; // @[LZD.scala 49:35]
  assign _T_164 = {_T_157,_T_159,_T_162}; // @[Cat.scala 29:58]
  assign _T_165 = _T_139[3:0]; // @[LZD.scala 44:32]
  assign _T_166 = _T_165[3:2]; // @[LZD.scala 43:32]
  assign _T_167 = _T_166 != 2'h0; // @[LZD.scala 39:14]
  assign _T_168 = _T_166[1]; // @[LZD.scala 39:21]
  assign _T_169 = _T_166[0]; // @[LZD.scala 39:30]
  assign _T_170 = ~ _T_169; // @[LZD.scala 39:27]
  assign _T_171 = _T_168 | _T_170; // @[LZD.scala 39:25]
  assign _T_172 = {_T_167,_T_171}; // @[Cat.scala 29:58]
  assign _T_173 = _T_165[1:0]; // @[LZD.scala 44:32]
  assign _T_174 = _T_173 != 2'h0; // @[LZD.scala 39:14]
  assign _T_175 = _T_173[1]; // @[LZD.scala 39:21]
  assign _T_176 = _T_173[0]; // @[LZD.scala 39:30]
  assign _T_177 = ~ _T_176; // @[LZD.scala 39:27]
  assign _T_178 = _T_175 | _T_177; // @[LZD.scala 39:25]
  assign _T_179 = {_T_174,_T_178}; // @[Cat.scala 29:58]
  assign _T_180 = _T_172[1]; // @[Shift.scala 12:21]
  assign _T_181 = _T_179[1]; // @[Shift.scala 12:21]
  assign _T_182 = _T_180 | _T_181; // @[LZD.scala 49:16]
  assign _T_183 = ~ _T_181; // @[LZD.scala 49:27]
  assign _T_184 = _T_180 | _T_183; // @[LZD.scala 49:25]
  assign _T_185 = _T_172[0:0]; // @[LZD.scala 49:47]
  assign _T_186 = _T_179[0:0]; // @[LZD.scala 49:59]
  assign _T_187 = _T_180 ? _T_185 : _T_186; // @[LZD.scala 49:35]
  assign _T_189 = {_T_182,_T_184,_T_187}; // @[Cat.scala 29:58]
  assign _T_190 = _T_164[2]; // @[Shift.scala 12:21]
  assign _T_191 = _T_189[2]; // @[Shift.scala 12:21]
  assign _T_192 = _T_190 | _T_191; // @[LZD.scala 49:16]
  assign _T_193 = ~ _T_191; // @[LZD.scala 49:27]
  assign _T_194 = _T_190 | _T_193; // @[LZD.scala 49:25]
  assign _T_195 = _T_164[1:0]; // @[LZD.scala 49:47]
  assign _T_196 = _T_189[1:0]; // @[LZD.scala 49:59]
  assign _T_197 = _T_190 ? _T_195 : _T_196; // @[LZD.scala 49:35]
  assign _T_199 = {_T_192,_T_194,_T_197}; // @[Cat.scala 29:58]
  assign _T_200 = _T_138[1:0]; // @[LZD.scala 44:32]
  assign _T_201 = _T_200 != 2'h0; // @[LZD.scala 39:14]
  assign _T_202 = _T_200[1]; // @[LZD.scala 39:21]
  assign _T_203 = _T_200[0]; // @[LZD.scala 39:30]
  assign _T_204 = ~ _T_203; // @[LZD.scala 39:27]
  assign _T_205 = _T_202 | _T_204; // @[LZD.scala 39:25]
  assign _T_207 = _T_199[3]; // @[Shift.scala 12:21]
  assign _T_209 = {1'h1,_T_201,_T_205}; // @[Cat.scala 29:58]
  assign _T_210 = _T_199[2:0]; // @[LZD.scala 55:32]
  assign _T_211 = _T_207 ? _T_210 : _T_209; // @[LZD.scala 55:20]
  assign _T_212 = {_T_207,_T_211}; // @[Cat.scala 29:58]
  assign _T_213 = ~ _T_212; // @[convert.scala 21:22]
  assign _T_214 = io_B[8:0]; // @[convert.scala 22:36]
  assign _T_215 = _T_213 < 4'h9; // @[Shift.scala 16:24]
  assign _T_217 = _T_213[3]; // @[Shift.scala 12:21]
  assign _T_218 = _T_214[0:0]; // @[Shift.scala 64:52]
  assign _T_220 = {_T_218,8'h0}; // @[Cat.scala 29:58]
  assign _T_221 = _T_217 ? _T_220 : _T_214; // @[Shift.scala 64:27]
  assign _T_222 = _T_213[2:0]; // @[Shift.scala 66:70]
  assign _T_223 = _T_222[2]; // @[Shift.scala 12:21]
  assign _T_224 = _T_221[4:0]; // @[Shift.scala 64:52]
  assign _T_226 = {_T_224,4'h0}; // @[Cat.scala 29:58]
  assign _T_227 = _T_223 ? _T_226 : _T_221; // @[Shift.scala 64:27]
  assign _T_228 = _T_222[1:0]; // @[Shift.scala 66:70]
  assign _T_229 = _T_228[1]; // @[Shift.scala 12:21]
  assign _T_230 = _T_227[6:0]; // @[Shift.scala 64:52]
  assign _T_232 = {_T_230,2'h0}; // @[Cat.scala 29:58]
  assign _T_233 = _T_229 ? _T_232 : _T_227; // @[Shift.scala 64:27]
  assign _T_234 = _T_228[0:0]; // @[Shift.scala 66:70]
  assign _T_236 = _T_233[7:0]; // @[Shift.scala 64:52]
  assign _T_237 = {_T_236,1'h0}; // @[Cat.scala 29:58]
  assign _T_238 = _T_234 ? _T_237 : _T_233; // @[Shift.scala 64:27]
  assign _T_239 = _T_215 ? _T_238 : 9'h0; // @[Shift.scala 16:10]
  assign _T_240 = _T_239[8:8]; // @[convert.scala 23:34]
  assign decB_fraction = _T_239[7:0]; // @[convert.scala 24:34]
  assign _T_242 = _T_135 == 1'h0; // @[convert.scala 25:26]
  assign _T_244 = _T_135 ? _T_213 : _T_212; // @[convert.scala 25:42]
  assign _T_247 = ~ _T_240; // @[convert.scala 26:67]
  assign _T_248 = _T_133 ? _T_247 : _T_240; // @[convert.scala 26:51]
  assign _T_249 = {_T_242,_T_244,_T_248}; // @[Cat.scala 29:58]
  assign _T_251 = io_B[10:0]; // @[convert.scala 29:56]
  assign _T_252 = _T_251 != 11'h0; // @[convert.scala 29:60]
  assign _T_253 = ~ _T_252; // @[convert.scala 29:41]
  assign decB_isNaR = _T_133 & _T_253; // @[convert.scala 29:39]
  assign _T_256 = _T_133 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_256 & _T_253; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_249); // @[convert.scala 32:24]
  assign aGTb = $signed(decA_scale) > $signed(decB_scale); // @[PositAdder.scala 24:32]
  assign greaterSign = aGTb ? _T_1 : _T_133; // @[PositAdder.scala 25:24]
  assign smallerSign = aGTb ? _T_133 : _T_1; // @[PositAdder.scala 26:24]
  assign greaterExp = aGTb ? $signed(decA_scale) : $signed(decB_scale); // @[PositAdder.scala 27:24]
  assign smallerExp = aGTb ? $signed(decB_scale) : $signed(decA_scale); // @[PositAdder.scala 28:24]
  assign greaterFrac = aGTb ? decA_fraction : decB_fraction; // @[PositAdder.scala 29:24]
  assign smallerFrac = aGTb ? decB_fraction : decA_fraction; // @[PositAdder.scala 30:24]
  assign smallerZero = aGTb ? decB_isZero : decA_isZero; // @[PositAdder.scala 31:24]
  assign _T_265 = $signed(greaterExp) - $signed(smallerExp); // @[PositAdder.scala 32:32]
  assign scale_diff = $signed(_T_265); // @[PositAdder.scala 32:32]
  assign _T_266 = ~ greaterSign; // @[PositAdder.scala 33:38]
  assign greaterSig = {greaterSign,_T_266,greaterFrac}; // @[Cat.scala 29:58]
  assign _T_268 = smallerSign | smallerZero; // @[PositAdder.scala 34:52]
  assign _T_269 = ~ _T_268; // @[PositAdder.scala 34:38]
  assign _T_272 = {smallerSign,_T_269,smallerFrac,3'h0}; // @[Cat.scala 29:58]
  assign _T_273 = $unsigned(scale_diff); // @[PositAdder.scala 35:68]
  assign _T_274 = _T_273 < 6'hd; // @[Shift.scala 39:24]
  assign _T_275 = _T_273[3:0]; // @[Shift.scala 40:44]
  assign _T_276 = _T_272[12:8]; // @[Shift.scala 90:30]
  assign _T_277 = _T_272[7:0]; // @[Shift.scala 90:48]
  assign _T_278 = _T_277 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_0 = {{4'd0}, _T_278}; // @[Shift.scala 90:39]
  assign _T_279 = _T_276 | _GEN_0; // @[Shift.scala 90:39]
  assign _T_280 = _T_275[3]; // @[Shift.scala 12:21]
  assign _T_281 = _T_272[12]; // @[Shift.scala 12:21]
  assign _T_283 = _T_281 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_284 = {_T_283,_T_279}; // @[Cat.scala 29:58]
  assign _T_285 = _T_280 ? _T_284 : _T_272; // @[Shift.scala 91:22]
  assign _T_286 = _T_275[2:0]; // @[Shift.scala 92:77]
  assign _T_287 = _T_285[12:4]; // @[Shift.scala 90:30]
  assign _T_288 = _T_285[3:0]; // @[Shift.scala 90:48]
  assign _T_289 = _T_288 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_1 = {{8'd0}, _T_289}; // @[Shift.scala 90:39]
  assign _T_290 = _T_287 | _GEN_1; // @[Shift.scala 90:39]
  assign _T_291 = _T_286[2]; // @[Shift.scala 12:21]
  assign _T_292 = _T_285[12]; // @[Shift.scala 12:21]
  assign _T_294 = _T_292 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_295 = {_T_294,_T_290}; // @[Cat.scala 29:58]
  assign _T_296 = _T_291 ? _T_295 : _T_285; // @[Shift.scala 91:22]
  assign _T_297 = _T_286[1:0]; // @[Shift.scala 92:77]
  assign _T_298 = _T_296[12:2]; // @[Shift.scala 90:30]
  assign _T_299 = _T_296[1:0]; // @[Shift.scala 90:48]
  assign _T_300 = _T_299 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_2 = {{10'd0}, _T_300}; // @[Shift.scala 90:39]
  assign _T_301 = _T_298 | _GEN_2; // @[Shift.scala 90:39]
  assign _T_302 = _T_297[1]; // @[Shift.scala 12:21]
  assign _T_303 = _T_296[12]; // @[Shift.scala 12:21]
  assign _T_305 = _T_303 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_306 = {_T_305,_T_301}; // @[Cat.scala 29:58]
  assign _T_307 = _T_302 ? _T_306 : _T_296; // @[Shift.scala 91:22]
  assign _T_308 = _T_297[0:0]; // @[Shift.scala 92:77]
  assign _T_309 = _T_307[12:1]; // @[Shift.scala 90:30]
  assign _T_310 = _T_307[0:0]; // @[Shift.scala 90:48]
  assign _GEN_3 = {{11'd0}, _T_310}; // @[Shift.scala 90:39]
  assign _T_312 = _T_309 | _GEN_3; // @[Shift.scala 90:39]
  assign _T_314 = _T_307[12]; // @[Shift.scala 12:21]
  assign _T_315 = {_T_314,_T_312}; // @[Cat.scala 29:58]
  assign _T_316 = _T_308 ? _T_315 : _T_307; // @[Shift.scala 91:22]
  assign _T_319 = _T_281 ? 13'h1fff : 13'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_274 ? _T_316 : _T_319; // @[Shift.scala 39:10]
  assign _T_320 = smallerSig[12:3]; // @[PositAdder.scala 36:45]
  assign rawSumSig = greaterSig + _T_320; // @[PositAdder.scala 36:32]
  assign _T_321 = _T_1 ^ _T_133; // @[PositAdder.scala 37:31]
  assign _T_322 = rawSumSig[10:10]; // @[PositAdder.scala 37:59]
  assign sumSign = _T_321 ^ _T_322; // @[PositAdder.scala 37:43]
  assign _T_323 = greaterSig + _T_320; // @[PositAdder.scala 38:48]
  assign _T_324 = smallerSig[2:0]; // @[PositAdder.scala 38:63]
  assign signSumSig = {sumSign,_T_323,_T_324}; // @[Cat.scala 29:58]
  assign _T_326 = signSumSig[13:1]; // @[PositAdder.scala 40:31]
  assign _T_327 = signSumSig[12:0]; // @[PositAdder.scala 40:66]
  assign sumXor = _T_326 ^ _T_327; // @[PositAdder.scala 40:49]
  assign _T_328 = sumXor[12:5]; // @[LZD.scala 43:32]
  assign _T_329 = _T_328[7:4]; // @[LZD.scala 43:32]
  assign _T_330 = _T_329[3:2]; // @[LZD.scala 43:32]
  assign _T_331 = _T_330 != 2'h0; // @[LZD.scala 39:14]
  assign _T_332 = _T_330[1]; // @[LZD.scala 39:21]
  assign _T_333 = _T_330[0]; // @[LZD.scala 39:30]
  assign _T_334 = ~ _T_333; // @[LZD.scala 39:27]
  assign _T_335 = _T_332 | _T_334; // @[LZD.scala 39:25]
  assign _T_336 = {_T_331,_T_335}; // @[Cat.scala 29:58]
  assign _T_337 = _T_329[1:0]; // @[LZD.scala 44:32]
  assign _T_338 = _T_337 != 2'h0; // @[LZD.scala 39:14]
  assign _T_339 = _T_337[1]; // @[LZD.scala 39:21]
  assign _T_340 = _T_337[0]; // @[LZD.scala 39:30]
  assign _T_341 = ~ _T_340; // @[LZD.scala 39:27]
  assign _T_342 = _T_339 | _T_341; // @[LZD.scala 39:25]
  assign _T_343 = {_T_338,_T_342}; // @[Cat.scala 29:58]
  assign _T_344 = _T_336[1]; // @[Shift.scala 12:21]
  assign _T_345 = _T_343[1]; // @[Shift.scala 12:21]
  assign _T_346 = _T_344 | _T_345; // @[LZD.scala 49:16]
  assign _T_347 = ~ _T_345; // @[LZD.scala 49:27]
  assign _T_348 = _T_344 | _T_347; // @[LZD.scala 49:25]
  assign _T_349 = _T_336[0:0]; // @[LZD.scala 49:47]
  assign _T_350 = _T_343[0:0]; // @[LZD.scala 49:59]
  assign _T_351 = _T_344 ? _T_349 : _T_350; // @[LZD.scala 49:35]
  assign _T_353 = {_T_346,_T_348,_T_351}; // @[Cat.scala 29:58]
  assign _T_354 = _T_328[3:0]; // @[LZD.scala 44:32]
  assign _T_355 = _T_354[3:2]; // @[LZD.scala 43:32]
  assign _T_356 = _T_355 != 2'h0; // @[LZD.scala 39:14]
  assign _T_357 = _T_355[1]; // @[LZD.scala 39:21]
  assign _T_358 = _T_355[0]; // @[LZD.scala 39:30]
  assign _T_359 = ~ _T_358; // @[LZD.scala 39:27]
  assign _T_360 = _T_357 | _T_359; // @[LZD.scala 39:25]
  assign _T_361 = {_T_356,_T_360}; // @[Cat.scala 29:58]
  assign _T_362 = _T_354[1:0]; // @[LZD.scala 44:32]
  assign _T_363 = _T_362 != 2'h0; // @[LZD.scala 39:14]
  assign _T_364 = _T_362[1]; // @[LZD.scala 39:21]
  assign _T_365 = _T_362[0]; // @[LZD.scala 39:30]
  assign _T_366 = ~ _T_365; // @[LZD.scala 39:27]
  assign _T_367 = _T_364 | _T_366; // @[LZD.scala 39:25]
  assign _T_368 = {_T_363,_T_367}; // @[Cat.scala 29:58]
  assign _T_369 = _T_361[1]; // @[Shift.scala 12:21]
  assign _T_370 = _T_368[1]; // @[Shift.scala 12:21]
  assign _T_371 = _T_369 | _T_370; // @[LZD.scala 49:16]
  assign _T_372 = ~ _T_370; // @[LZD.scala 49:27]
  assign _T_373 = _T_369 | _T_372; // @[LZD.scala 49:25]
  assign _T_374 = _T_361[0:0]; // @[LZD.scala 49:47]
  assign _T_375 = _T_368[0:0]; // @[LZD.scala 49:59]
  assign _T_376 = _T_369 ? _T_374 : _T_375; // @[LZD.scala 49:35]
  assign _T_378 = {_T_371,_T_373,_T_376}; // @[Cat.scala 29:58]
  assign _T_379 = _T_353[2]; // @[Shift.scala 12:21]
  assign _T_380 = _T_378[2]; // @[Shift.scala 12:21]
  assign _T_381 = _T_379 | _T_380; // @[LZD.scala 49:16]
  assign _T_382 = ~ _T_380; // @[LZD.scala 49:27]
  assign _T_383 = _T_379 | _T_382; // @[LZD.scala 49:25]
  assign _T_384 = _T_353[1:0]; // @[LZD.scala 49:47]
  assign _T_385 = _T_378[1:0]; // @[LZD.scala 49:59]
  assign _T_386 = _T_379 ? _T_384 : _T_385; // @[LZD.scala 49:35]
  assign _T_388 = {_T_381,_T_383,_T_386}; // @[Cat.scala 29:58]
  assign _T_389 = sumXor[4:0]; // @[LZD.scala 44:32]
  assign _T_390 = _T_389[4:1]; // @[LZD.scala 43:32]
  assign _T_391 = _T_390[3:2]; // @[LZD.scala 43:32]
  assign _T_392 = _T_391 != 2'h0; // @[LZD.scala 39:14]
  assign _T_393 = _T_391[1]; // @[LZD.scala 39:21]
  assign _T_394 = _T_391[0]; // @[LZD.scala 39:30]
  assign _T_395 = ~ _T_394; // @[LZD.scala 39:27]
  assign _T_396 = _T_393 | _T_395; // @[LZD.scala 39:25]
  assign _T_397 = {_T_392,_T_396}; // @[Cat.scala 29:58]
  assign _T_398 = _T_390[1:0]; // @[LZD.scala 44:32]
  assign _T_399 = _T_398 != 2'h0; // @[LZD.scala 39:14]
  assign _T_400 = _T_398[1]; // @[LZD.scala 39:21]
  assign _T_401 = _T_398[0]; // @[LZD.scala 39:30]
  assign _T_402 = ~ _T_401; // @[LZD.scala 39:27]
  assign _T_403 = _T_400 | _T_402; // @[LZD.scala 39:25]
  assign _T_404 = {_T_399,_T_403}; // @[Cat.scala 29:58]
  assign _T_405 = _T_397[1]; // @[Shift.scala 12:21]
  assign _T_406 = _T_404[1]; // @[Shift.scala 12:21]
  assign _T_407 = _T_405 | _T_406; // @[LZD.scala 49:16]
  assign _T_408 = ~ _T_406; // @[LZD.scala 49:27]
  assign _T_409 = _T_405 | _T_408; // @[LZD.scala 49:25]
  assign _T_410 = _T_397[0:0]; // @[LZD.scala 49:47]
  assign _T_411 = _T_404[0:0]; // @[LZD.scala 49:59]
  assign _T_412 = _T_405 ? _T_410 : _T_411; // @[LZD.scala 49:35]
  assign _T_414 = {_T_407,_T_409,_T_412}; // @[Cat.scala 29:58]
  assign _T_415 = _T_389[0:0]; // @[LZD.scala 44:32]
  assign _T_417 = _T_414[2]; // @[Shift.scala 12:21]
  assign _T_419 = {1'h1,_T_415}; // @[Cat.scala 29:58]
  assign _T_420 = _T_414[1:0]; // @[LZD.scala 55:32]
  assign _T_421 = _T_417 ? _T_420 : _T_419; // @[LZD.scala 55:20]
  assign _T_422 = {_T_417,_T_421}; // @[Cat.scala 29:58]
  assign _T_423 = _T_388[3]; // @[Shift.scala 12:21]
  assign _T_425 = _T_388[2:0]; // @[LZD.scala 55:32]
  assign _T_426 = _T_423 ? _T_425 : _T_422; // @[LZD.scala 55:20]
  assign sumLZD = {_T_423,_T_426}; // @[Cat.scala 29:58]
  assign _T_427 = {1'h1,_T_423,_T_426}; // @[Cat.scala 29:58]
  assign _T_428 = $signed(_T_427); // @[PositAdder.scala 42:38]
  assign _T_430 = $signed(_T_428) + $signed(5'sh2); // @[PositAdder.scala 42:45]
  assign scaleBias = $signed(_T_430); // @[PositAdder.scala 42:45]
  assign _GEN_4 = {{1{scaleBias[4]}},scaleBias}; // @[PositAdder.scala 43:32]
  assign sumScale = $signed(greaterExp) + $signed(_GEN_4); // @[PositAdder.scala 43:32]
  assign overflow = $signed(sumScale) > $signed(7'sh14); // @[PositAdder.scala 44:30]
  assign normalShift = ~ sumLZD; // @[PositAdder.scala 45:22]
  assign _T_431 = signSumSig[11:0]; // @[PositAdder.scala 46:36]
  assign _T_432 = normalShift < 4'hc; // @[Shift.scala 16:24]
  assign _T_434 = normalShift[3]; // @[Shift.scala 12:21]
  assign _T_435 = _T_431[3:0]; // @[Shift.scala 64:52]
  assign _T_437 = {_T_435,8'h0}; // @[Cat.scala 29:58]
  assign _T_438 = _T_434 ? _T_437 : _T_431; // @[Shift.scala 64:27]
  assign _T_439 = normalShift[2:0]; // @[Shift.scala 66:70]
  assign _T_440 = _T_439[2]; // @[Shift.scala 12:21]
  assign _T_441 = _T_438[7:0]; // @[Shift.scala 64:52]
  assign _T_443 = {_T_441,4'h0}; // @[Cat.scala 29:58]
  assign _T_444 = _T_440 ? _T_443 : _T_438; // @[Shift.scala 64:27]
  assign _T_445 = _T_439[1:0]; // @[Shift.scala 66:70]
  assign _T_446 = _T_445[1]; // @[Shift.scala 12:21]
  assign _T_447 = _T_444[9:0]; // @[Shift.scala 64:52]
  assign _T_449 = {_T_447,2'h0}; // @[Cat.scala 29:58]
  assign _T_450 = _T_446 ? _T_449 : _T_444; // @[Shift.scala 64:27]
  assign _T_451 = _T_445[0:0]; // @[Shift.scala 66:70]
  assign _T_453 = _T_450[10:0]; // @[Shift.scala 64:52]
  assign _T_454 = {_T_453,1'h0}; // @[Cat.scala 29:58]
  assign _T_455 = _T_451 ? _T_454 : _T_450; // @[Shift.scala 64:27]
  assign shiftSig = _T_432 ? _T_455 : 12'h0; // @[Shift.scala 16:10]
  assign _T_456 = overflow ? $signed(7'sh14) : $signed(sumScale); // @[PositAdder.scala 51:24]
  assign decS_fraction = shiftSig[11:4]; // @[PositAdder.scala 52:34]
  assign decS_isNaR = decA_isNaR | decB_isNaR; // @[PositAdder.scala 53:32]
  assign _T_459 = signSumSig != 14'h0; // @[PositAdder.scala 54:33]
  assign _T_460 = ~ _T_459; // @[PositAdder.scala 54:21]
  assign _T_461 = decA_isZero & decB_isZero; // @[PositAdder.scala 54:52]
  assign decS_isZero = _T_460 | _T_461; // @[PositAdder.scala 54:37]
  assign _T_463 = shiftSig[3:2]; // @[PositAdder.scala 55:33]
  assign _T_464 = shiftSig[1]; // @[PositAdder.scala 55:49]
  assign _T_465 = shiftSig[0]; // @[PositAdder.scala 55:63]
  assign _T_466 = _T_464 | _T_465; // @[PositAdder.scala 55:53]
  assign _GEN_5 = _T_456[5:0]; // @[PositAdder.scala 48:25 PositAdder.scala 51:18]
  assign decS_scale = $signed(_GEN_5); // @[PositAdder.scala 48:25 PositAdder.scala 51:18]
  assign _T_469 = decS_scale[0]; // @[convert.scala 46:61]
  assign _T_470 = ~ _T_469; // @[convert.scala 46:52]
  assign _T_472 = sumSign ? _T_470 : _T_469; // @[convert.scala 46:42]
  assign _T_473 = decS_scale[5:1]; // @[convert.scala 48:34]
  assign _T_474 = _T_473[4:4]; // @[convert.scala 49:36]
  assign _T_476 = ~ _T_473; // @[convert.scala 50:36]
  assign _T_477 = $signed(_T_476); // @[convert.scala 50:36]
  assign _T_478 = _T_474 ? $signed(_T_477) : $signed(_T_473); // @[convert.scala 50:28]
  assign _T_479 = _T_474 ^ sumSign; // @[convert.scala 51:31]
  assign _T_480 = ~ _T_479; // @[convert.scala 52:43]
  assign _T_484 = {_T_480,_T_479,_T_472,decS_fraction,_T_463,_T_466}; // @[Cat.scala 29:58]
  assign _T_485 = $unsigned(_T_478); // @[Shift.scala 39:17]
  assign _T_486 = _T_485 < 5'he; // @[Shift.scala 39:24]
  assign _T_487 = _T_478[3:0]; // @[Shift.scala 40:44]
  assign _T_488 = _T_484[13:8]; // @[Shift.scala 90:30]
  assign _T_489 = _T_484[7:0]; // @[Shift.scala 90:48]
  assign _T_490 = _T_489 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_6 = {{5'd0}, _T_490}; // @[Shift.scala 90:39]
  assign _T_491 = _T_488 | _GEN_6; // @[Shift.scala 90:39]
  assign _T_492 = _T_487[3]; // @[Shift.scala 12:21]
  assign _T_493 = _T_484[13]; // @[Shift.scala 12:21]
  assign _T_495 = _T_493 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_496 = {_T_495,_T_491}; // @[Cat.scala 29:58]
  assign _T_497 = _T_492 ? _T_496 : _T_484; // @[Shift.scala 91:22]
  assign _T_498 = _T_487[2:0]; // @[Shift.scala 92:77]
  assign _T_499 = _T_497[13:4]; // @[Shift.scala 90:30]
  assign _T_500 = _T_497[3:0]; // @[Shift.scala 90:48]
  assign _T_501 = _T_500 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_7 = {{9'd0}, _T_501}; // @[Shift.scala 90:39]
  assign _T_502 = _T_499 | _GEN_7; // @[Shift.scala 90:39]
  assign _T_503 = _T_498[2]; // @[Shift.scala 12:21]
  assign _T_504 = _T_497[13]; // @[Shift.scala 12:21]
  assign _T_506 = _T_504 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_507 = {_T_506,_T_502}; // @[Cat.scala 29:58]
  assign _T_508 = _T_503 ? _T_507 : _T_497; // @[Shift.scala 91:22]
  assign _T_509 = _T_498[1:0]; // @[Shift.scala 92:77]
  assign _T_510 = _T_508[13:2]; // @[Shift.scala 90:30]
  assign _T_511 = _T_508[1:0]; // @[Shift.scala 90:48]
  assign _T_512 = _T_511 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_8 = {{11'd0}, _T_512}; // @[Shift.scala 90:39]
  assign _T_513 = _T_510 | _GEN_8; // @[Shift.scala 90:39]
  assign _T_514 = _T_509[1]; // @[Shift.scala 12:21]
  assign _T_515 = _T_508[13]; // @[Shift.scala 12:21]
  assign _T_517 = _T_515 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_518 = {_T_517,_T_513}; // @[Cat.scala 29:58]
  assign _T_519 = _T_514 ? _T_518 : _T_508; // @[Shift.scala 91:22]
  assign _T_520 = _T_509[0:0]; // @[Shift.scala 92:77]
  assign _T_521 = _T_519[13:1]; // @[Shift.scala 90:30]
  assign _T_522 = _T_519[0:0]; // @[Shift.scala 90:48]
  assign _GEN_9 = {{12'd0}, _T_522}; // @[Shift.scala 90:39]
  assign _T_524 = _T_521 | _GEN_9; // @[Shift.scala 90:39]
  assign _T_526 = _T_519[13]; // @[Shift.scala 12:21]
  assign _T_527 = {_T_526,_T_524}; // @[Cat.scala 29:58]
  assign _T_528 = _T_520 ? _T_527 : _T_519; // @[Shift.scala 91:22]
  assign _T_531 = _T_493 ? 14'h3fff : 14'h0; // @[Bitwise.scala 71:12]
  assign _T_532 = _T_486 ? _T_528 : _T_531; // @[Shift.scala 39:10]
  assign _T_533 = _T_532[3]; // @[convert.scala 55:31]
  assign _T_534 = _T_532[2]; // @[convert.scala 56:31]
  assign _T_535 = _T_532[1]; // @[convert.scala 57:31]
  assign _T_536 = _T_532[0]; // @[convert.scala 58:31]
  assign _T_537 = _T_532[13:3]; // @[convert.scala 59:69]
  assign _T_538 = _T_537 != 11'h0; // @[convert.scala 59:81]
  assign _T_539 = ~ _T_538; // @[convert.scala 59:50]
  assign _T_541 = _T_537 == 11'h7ff; // @[convert.scala 60:81]
  assign _T_542 = _T_533 | _T_535; // @[convert.scala 61:44]
  assign _T_543 = _T_542 | _T_536; // @[convert.scala 61:52]
  assign _T_544 = _T_534 & _T_543; // @[convert.scala 61:36]
  assign _T_545 = ~ _T_541; // @[convert.scala 62:63]
  assign _T_546 = _T_545 & _T_544; // @[convert.scala 62:103]
  assign _T_547 = _T_539 | _T_546; // @[convert.scala 62:60]
  assign _GEN_10 = {{10'd0}, _T_547}; // @[convert.scala 63:56]
  assign _T_550 = _T_537 + _GEN_10; // @[convert.scala 63:56]
  assign _T_551 = {sumSign,_T_550}; // @[Cat.scala 29:58]
  assign _T_553 = decS_isZero ? 12'h0 : _T_551; // @[Mux.scala 87:16]
  assign io_S = decS_isNaR ? 12'h800 : _T_553; // @[PositAdder.scala 57:8]
endmodule
