module PositMultiplier8_1(
  input        clock,
  input        reset,
  input  [7:0] io_A,
  input  [7:0] io_B,
  output [7:0] io_M
);
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [5:0] _T_4; // @[convert.scala 19:24]
  wire [5:0] _T_5; // @[convert.scala 19:43]
  wire [5:0] _T_6; // @[convert.scala 19:39]
  wire [3:0] _T_7; // @[LZD.scala 43:32]
  wire [1:0] _T_8; // @[LZD.scala 43:32]
  wire  _T_9; // @[LZD.scala 39:14]
  wire  _T_10; // @[LZD.scala 39:21]
  wire  _T_11; // @[LZD.scala 39:30]
  wire  _T_12; // @[LZD.scala 39:27]
  wire  _T_13; // @[LZD.scala 39:25]
  wire [1:0] _T_14; // @[Cat.scala 29:58]
  wire [1:0] _T_15; // @[LZD.scala 44:32]
  wire  _T_16; // @[LZD.scala 39:14]
  wire  _T_17; // @[LZD.scala 39:21]
  wire  _T_18; // @[LZD.scala 39:30]
  wire  _T_19; // @[LZD.scala 39:27]
  wire  _T_20; // @[LZD.scala 39:25]
  wire [1:0] _T_21; // @[Cat.scala 29:58]
  wire  _T_22; // @[Shift.scala 12:21]
  wire  _T_23; // @[Shift.scala 12:21]
  wire  _T_24; // @[LZD.scala 49:16]
  wire  _T_25; // @[LZD.scala 49:27]
  wire  _T_26; // @[LZD.scala 49:25]
  wire  _T_27; // @[LZD.scala 49:47]
  wire  _T_28; // @[LZD.scala 49:59]
  wire  _T_29; // @[LZD.scala 49:35]
  wire [2:0] _T_31; // @[Cat.scala 29:58]
  wire [1:0] _T_32; // @[LZD.scala 44:32]
  wire  _T_33; // @[LZD.scala 39:14]
  wire  _T_34; // @[LZD.scala 39:21]
  wire  _T_35; // @[LZD.scala 39:30]
  wire  _T_36; // @[LZD.scala 39:27]
  wire  _T_37; // @[LZD.scala 39:25]
  wire [1:0] _T_38; // @[Cat.scala 29:58]
  wire  _T_39; // @[Shift.scala 12:21]
  wire [1:0] _T_41; // @[LZD.scala 55:32]
  wire [1:0] _T_42; // @[LZD.scala 55:20]
  wire [2:0] _T_43; // @[Cat.scala 29:58]
  wire [2:0] _T_44; // @[convert.scala 21:22]
  wire [4:0] _T_45; // @[convert.scala 22:36]
  wire  _T_46; // @[Shift.scala 16:24]
  wire  _T_48; // @[Shift.scala 12:21]
  wire  _T_49; // @[Shift.scala 64:52]
  wire [4:0] _T_51; // @[Cat.scala 29:58]
  wire [4:0] _T_52; // @[Shift.scala 64:27]
  wire [1:0] _T_53; // @[Shift.scala 66:70]
  wire  _T_54; // @[Shift.scala 12:21]
  wire [2:0] _T_55; // @[Shift.scala 64:52]
  wire [4:0] _T_57; // @[Cat.scala 29:58]
  wire [4:0] _T_58; // @[Shift.scala 64:27]
  wire  _T_59; // @[Shift.scala 66:70]
  wire [3:0] _T_61; // @[Shift.scala 64:52]
  wire [4:0] _T_62; // @[Cat.scala 29:58]
  wire [4:0] _T_63; // @[Shift.scala 64:27]
  wire [4:0] _T_64; // @[Shift.scala 16:10]
  wire  _T_65; // @[convert.scala 23:34]
  wire [3:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_67; // @[convert.scala 25:26]
  wire [2:0] _T_69; // @[convert.scala 25:42]
  wire  _T_72; // @[convert.scala 26:67]
  wire  _T_73; // @[convert.scala 26:51]
  wire [4:0] _T_74; // @[Cat.scala 29:58]
  wire [6:0] _T_76; // @[convert.scala 29:56]
  wire  _T_77; // @[convert.scala 29:60]
  wire  _T_78; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_81; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [4:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_90; // @[convert.scala 18:24]
  wire  _T_91; // @[convert.scala 18:40]
  wire  _T_92; // @[convert.scala 18:36]
  wire [5:0] _T_93; // @[convert.scala 19:24]
  wire [5:0] _T_94; // @[convert.scala 19:43]
  wire [5:0] _T_95; // @[convert.scala 19:39]
  wire [3:0] _T_96; // @[LZD.scala 43:32]
  wire [1:0] _T_97; // @[LZD.scala 43:32]
  wire  _T_98; // @[LZD.scala 39:14]
  wire  _T_99; // @[LZD.scala 39:21]
  wire  _T_100; // @[LZD.scala 39:30]
  wire  _T_101; // @[LZD.scala 39:27]
  wire  _T_102; // @[LZD.scala 39:25]
  wire [1:0] _T_103; // @[Cat.scala 29:58]
  wire [1:0] _T_104; // @[LZD.scala 44:32]
  wire  _T_105; // @[LZD.scala 39:14]
  wire  _T_106; // @[LZD.scala 39:21]
  wire  _T_107; // @[LZD.scala 39:30]
  wire  _T_108; // @[LZD.scala 39:27]
  wire  _T_109; // @[LZD.scala 39:25]
  wire [1:0] _T_110; // @[Cat.scala 29:58]
  wire  _T_111; // @[Shift.scala 12:21]
  wire  _T_112; // @[Shift.scala 12:21]
  wire  _T_113; // @[LZD.scala 49:16]
  wire  _T_114; // @[LZD.scala 49:27]
  wire  _T_115; // @[LZD.scala 49:25]
  wire  _T_116; // @[LZD.scala 49:47]
  wire  _T_117; // @[LZD.scala 49:59]
  wire  _T_118; // @[LZD.scala 49:35]
  wire [2:0] _T_120; // @[Cat.scala 29:58]
  wire [1:0] _T_121; // @[LZD.scala 44:32]
  wire  _T_122; // @[LZD.scala 39:14]
  wire  _T_123; // @[LZD.scala 39:21]
  wire  _T_124; // @[LZD.scala 39:30]
  wire  _T_125; // @[LZD.scala 39:27]
  wire  _T_126; // @[LZD.scala 39:25]
  wire [1:0] _T_127; // @[Cat.scala 29:58]
  wire  _T_128; // @[Shift.scala 12:21]
  wire [1:0] _T_130; // @[LZD.scala 55:32]
  wire [1:0] _T_131; // @[LZD.scala 55:20]
  wire [2:0] _T_132; // @[Cat.scala 29:58]
  wire [2:0] _T_133; // @[convert.scala 21:22]
  wire [4:0] _T_134; // @[convert.scala 22:36]
  wire  _T_135; // @[Shift.scala 16:24]
  wire  _T_137; // @[Shift.scala 12:21]
  wire  _T_138; // @[Shift.scala 64:52]
  wire [4:0] _T_140; // @[Cat.scala 29:58]
  wire [4:0] _T_141; // @[Shift.scala 64:27]
  wire [1:0] _T_142; // @[Shift.scala 66:70]
  wire  _T_143; // @[Shift.scala 12:21]
  wire [2:0] _T_144; // @[Shift.scala 64:52]
  wire [4:0] _T_146; // @[Cat.scala 29:58]
  wire [4:0] _T_147; // @[Shift.scala 64:27]
  wire  _T_148; // @[Shift.scala 66:70]
  wire [3:0] _T_150; // @[Shift.scala 64:52]
  wire [4:0] _T_151; // @[Cat.scala 29:58]
  wire [4:0] _T_152; // @[Shift.scala 64:27]
  wire [4:0] _T_153; // @[Shift.scala 16:10]
  wire  _T_154; // @[convert.scala 23:34]
  wire [3:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_156; // @[convert.scala 25:26]
  wire [2:0] _T_158; // @[convert.scala 25:42]
  wire  _T_161; // @[convert.scala 26:67]
  wire  _T_162; // @[convert.scala 26:51]
  wire [4:0] _T_163; // @[Cat.scala 29:58]
  wire [6:0] _T_165; // @[convert.scala 29:56]
  wire  _T_166; // @[convert.scala 29:60]
  wire  _T_167; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_170; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [4:0] decB_scale; // @[convert.scala 32:24]
  wire  _T_178; // @[PositMultiplier.scala 43:34]
  wire [5:0] _T_180; // @[Cat.scala 29:58]
  wire [5:0] sigA; // @[PositMultiplier.scala 43:61]
  wire  _T_181; // @[PositMultiplier.scala 44:34]
  wire [5:0] _T_183; // @[Cat.scala 29:58]
  wire [5:0] sigB; // @[PositMultiplier.scala 44:61]
  wire [11:0] _T_184; // @[PositMultiplier.scala 45:25]
  wire [11:0] sigP; // @[PositMultiplier.scala 45:33]
  wire [1:0] head2; // @[PositMultiplier.scala 46:28]
  wire  _T_185; // @[PositMultiplier.scala 47:31]
  wire  _T_186; // @[PositMultiplier.scala 47:25]
  wire  _T_187; // @[PositMultiplier.scala 47:42]
  wire  addTwo; // @[PositMultiplier.scala 47:35]
  wire  _T_188; // @[PositMultiplier.scala 49:23]
  wire  _T_189; // @[PositMultiplier.scala 49:49]
  wire  addOne; // @[PositMultiplier.scala 49:43]
  wire [1:0] _T_190; // @[Cat.scala 29:58]
  wire [2:0] expBias; // @[PositMultiplier.scala 50:39]
  wire [8:0] _T_191; // @[PositMultiplier.scala 53:81]
  wire [7:0] _T_192; // @[PositMultiplier.scala 54:81]
  wire [8:0] _T_193; // @[PositMultiplier.scala 54:104]
  wire [8:0] frac; // @[PositMultiplier.scala 51:22]
  wire [5:0] _T_194; // @[PositMultiplier.scala 56:30]
  wire [5:0] _GEN_0; // @[PositMultiplier.scala 56:44]
  wire [5:0] _T_196; // @[PositMultiplier.scala 56:44]
  wire [5:0] mulScale; // @[PositMultiplier.scala 56:44]
  wire  underflow; // @[PositMultiplier.scala 57:28]
  wire  overflow; // @[PositMultiplier.scala 58:28]
  wire  decM_sign; // @[PositMultiplier.scala 62:29]
  wire [5:0] _T_199; // @[Mux.scala 87:16]
  wire [5:0] _T_200; // @[Mux.scala 87:16]
  wire [3:0] decM_fraction; // @[PositMultiplier.scala 70:29]
  wire  decM_isNaR; // @[PositMultiplier.scala 71:31]
  wire  decM_isZero; // @[PositMultiplier.scala 72:32]
  wire [4:0] grsTmp; // @[PositMultiplier.scala 75:30]
  wire [1:0] _T_204; // @[PositMultiplier.scala 78:32]
  wire [2:0] _T_205; // @[PositMultiplier.scala 78:48]
  wire  _T_206; // @[PositMultiplier.scala 78:52]
  wire [4:0] _GEN_1; // @[PositMultiplier.scala 60:23 PositMultiplier.scala 63:17]
  wire [4:0] decM_scale; // @[PositMultiplier.scala 60:23 PositMultiplier.scala 63:17]
  wire  _T_209; // @[convert.scala 46:61]
  wire  _T_210; // @[convert.scala 46:52]
  wire  _T_212; // @[convert.scala 46:42]
  wire [3:0] _T_213; // @[convert.scala 48:34]
  wire  _T_214; // @[convert.scala 49:36]
  wire [3:0] _T_216; // @[convert.scala 50:36]
  wire [3:0] _T_217; // @[convert.scala 50:36]
  wire [3:0] _T_218; // @[convert.scala 50:28]
  wire  _T_219; // @[convert.scala 51:31]
  wire  _T_220; // @[convert.scala 52:43]
  wire [9:0] _T_224; // @[Cat.scala 29:58]
  wire [3:0] _T_225; // @[Shift.scala 39:17]
  wire  _T_226; // @[Shift.scala 39:24]
  wire [1:0] _T_228; // @[Shift.scala 90:30]
  wire [7:0] _T_229; // @[Shift.scala 90:48]
  wire  _T_230; // @[Shift.scala 90:57]
  wire [1:0] _GEN_2; // @[Shift.scala 90:39]
  wire [1:0] _T_231; // @[Shift.scala 90:39]
  wire  _T_232; // @[Shift.scala 12:21]
  wire  _T_233; // @[Shift.scala 12:21]
  wire [7:0] _T_235; // @[Bitwise.scala 71:12]
  wire [9:0] _T_236; // @[Cat.scala 29:58]
  wire [9:0] _T_237; // @[Shift.scala 91:22]
  wire [2:0] _T_238; // @[Shift.scala 92:77]
  wire [5:0] _T_239; // @[Shift.scala 90:30]
  wire [3:0] _T_240; // @[Shift.scala 90:48]
  wire  _T_241; // @[Shift.scala 90:57]
  wire [5:0] _GEN_3; // @[Shift.scala 90:39]
  wire [5:0] _T_242; // @[Shift.scala 90:39]
  wire  _T_243; // @[Shift.scala 12:21]
  wire  _T_244; // @[Shift.scala 12:21]
  wire [3:0] _T_246; // @[Bitwise.scala 71:12]
  wire [9:0] _T_247; // @[Cat.scala 29:58]
  wire [9:0] _T_248; // @[Shift.scala 91:22]
  wire [1:0] _T_249; // @[Shift.scala 92:77]
  wire [7:0] _T_250; // @[Shift.scala 90:30]
  wire [1:0] _T_251; // @[Shift.scala 90:48]
  wire  _T_252; // @[Shift.scala 90:57]
  wire [7:0] _GEN_4; // @[Shift.scala 90:39]
  wire [7:0] _T_253; // @[Shift.scala 90:39]
  wire  _T_254; // @[Shift.scala 12:21]
  wire  _T_255; // @[Shift.scala 12:21]
  wire [1:0] _T_257; // @[Bitwise.scala 71:12]
  wire [9:0] _T_258; // @[Cat.scala 29:58]
  wire [9:0] _T_259; // @[Shift.scala 91:22]
  wire  _T_260; // @[Shift.scala 92:77]
  wire [8:0] _T_261; // @[Shift.scala 90:30]
  wire  _T_262; // @[Shift.scala 90:48]
  wire [8:0] _GEN_5; // @[Shift.scala 90:39]
  wire [8:0] _T_264; // @[Shift.scala 90:39]
  wire  _T_266; // @[Shift.scala 12:21]
  wire [9:0] _T_267; // @[Cat.scala 29:58]
  wire [9:0] _T_268; // @[Shift.scala 91:22]
  wire [9:0] _T_271; // @[Bitwise.scala 71:12]
  wire [9:0] _T_272; // @[Shift.scala 39:10]
  wire  _T_273; // @[convert.scala 55:31]
  wire  _T_274; // @[convert.scala 56:31]
  wire  _T_275; // @[convert.scala 57:31]
  wire  _T_276; // @[convert.scala 58:31]
  wire [6:0] _T_277; // @[convert.scala 59:69]
  wire  _T_278; // @[convert.scala 59:81]
  wire  _T_279; // @[convert.scala 59:50]
  wire  _T_281; // @[convert.scala 60:81]
  wire  _T_282; // @[convert.scala 61:44]
  wire  _T_283; // @[convert.scala 61:52]
  wire  _T_284; // @[convert.scala 61:36]
  wire  _T_285; // @[convert.scala 62:63]
  wire  _T_286; // @[convert.scala 62:103]
  wire  _T_287; // @[convert.scala 62:60]
  wire [6:0] _GEN_6; // @[convert.scala 63:56]
  wire [6:0] _T_290; // @[convert.scala 63:56]
  wire [7:0] _T_291; // @[Cat.scala 29:58]
  wire [7:0] _T_293; // @[Mux.scala 87:16]
  assign _T_1 = io_A[7]; // @[convert.scala 18:24]
  assign _T_2 = io_A[6]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[6:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[5:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[5:2]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[3:2]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8 != 2'h0; // @[LZD.scala 39:14]
  assign _T_10 = _T_8[1]; // @[LZD.scala 39:21]
  assign _T_11 = _T_8[0]; // @[LZD.scala 39:30]
  assign _T_12 = ~ _T_11; // @[LZD.scala 39:27]
  assign _T_13 = _T_10 | _T_12; // @[LZD.scala 39:25]
  assign _T_14 = {_T_9,_T_13}; // @[Cat.scala 29:58]
  assign _T_15 = _T_7[1:0]; // @[LZD.scala 44:32]
  assign _T_16 = _T_15 != 2'h0; // @[LZD.scala 39:14]
  assign _T_17 = _T_15[1]; // @[LZD.scala 39:21]
  assign _T_18 = _T_15[0]; // @[LZD.scala 39:30]
  assign _T_19 = ~ _T_18; // @[LZD.scala 39:27]
  assign _T_20 = _T_17 | _T_19; // @[LZD.scala 39:25]
  assign _T_21 = {_T_16,_T_20}; // @[Cat.scala 29:58]
  assign _T_22 = _T_14[1]; // @[Shift.scala 12:21]
  assign _T_23 = _T_21[1]; // @[Shift.scala 12:21]
  assign _T_24 = _T_22 | _T_23; // @[LZD.scala 49:16]
  assign _T_25 = ~ _T_23; // @[LZD.scala 49:27]
  assign _T_26 = _T_22 | _T_25; // @[LZD.scala 49:25]
  assign _T_27 = _T_14[0:0]; // @[LZD.scala 49:47]
  assign _T_28 = _T_21[0:0]; // @[LZD.scala 49:59]
  assign _T_29 = _T_22 ? _T_27 : _T_28; // @[LZD.scala 49:35]
  assign _T_31 = {_T_24,_T_26,_T_29}; // @[Cat.scala 29:58]
  assign _T_32 = _T_6[1:0]; // @[LZD.scala 44:32]
  assign _T_33 = _T_32 != 2'h0; // @[LZD.scala 39:14]
  assign _T_34 = _T_32[1]; // @[LZD.scala 39:21]
  assign _T_35 = _T_32[0]; // @[LZD.scala 39:30]
  assign _T_36 = ~ _T_35; // @[LZD.scala 39:27]
  assign _T_37 = _T_34 | _T_36; // @[LZD.scala 39:25]
  assign _T_38 = {_T_33,_T_37}; // @[Cat.scala 29:58]
  assign _T_39 = _T_31[2]; // @[Shift.scala 12:21]
  assign _T_41 = _T_31[1:0]; // @[LZD.scala 55:32]
  assign _T_42 = _T_39 ? _T_41 : _T_38; // @[LZD.scala 55:20]
  assign _T_43 = {_T_39,_T_42}; // @[Cat.scala 29:58]
  assign _T_44 = ~ _T_43; // @[convert.scala 21:22]
  assign _T_45 = io_A[4:0]; // @[convert.scala 22:36]
  assign _T_46 = _T_44 < 3'h5; // @[Shift.scala 16:24]
  assign _T_48 = _T_44[2]; // @[Shift.scala 12:21]
  assign _T_49 = _T_45[0:0]; // @[Shift.scala 64:52]
  assign _T_51 = {_T_49,4'h0}; // @[Cat.scala 29:58]
  assign _T_52 = _T_48 ? _T_51 : _T_45; // @[Shift.scala 64:27]
  assign _T_53 = _T_44[1:0]; // @[Shift.scala 66:70]
  assign _T_54 = _T_53[1]; // @[Shift.scala 12:21]
  assign _T_55 = _T_52[2:0]; // @[Shift.scala 64:52]
  assign _T_57 = {_T_55,2'h0}; // @[Cat.scala 29:58]
  assign _T_58 = _T_54 ? _T_57 : _T_52; // @[Shift.scala 64:27]
  assign _T_59 = _T_53[0:0]; // @[Shift.scala 66:70]
  assign _T_61 = _T_58[3:0]; // @[Shift.scala 64:52]
  assign _T_62 = {_T_61,1'h0}; // @[Cat.scala 29:58]
  assign _T_63 = _T_59 ? _T_62 : _T_58; // @[Shift.scala 64:27]
  assign _T_64 = _T_46 ? _T_63 : 5'h0; // @[Shift.scala 16:10]
  assign _T_65 = _T_64[4:4]; // @[convert.scala 23:34]
  assign decA_fraction = _T_64[3:0]; // @[convert.scala 24:34]
  assign _T_67 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_69 = _T_3 ? _T_44 : _T_43; // @[convert.scala 25:42]
  assign _T_72 = ~ _T_65; // @[convert.scala 26:67]
  assign _T_73 = _T_1 ? _T_72 : _T_65; // @[convert.scala 26:51]
  assign _T_74 = {_T_67,_T_69,_T_73}; // @[Cat.scala 29:58]
  assign _T_76 = io_A[6:0]; // @[convert.scala 29:56]
  assign _T_77 = _T_76 != 7'h0; // @[convert.scala 29:60]
  assign _T_78 = ~ _T_77; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_78; // @[convert.scala 29:39]
  assign _T_81 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_81 & _T_78; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_74); // @[convert.scala 32:24]
  assign _T_90 = io_B[7]; // @[convert.scala 18:24]
  assign _T_91 = io_B[6]; // @[convert.scala 18:40]
  assign _T_92 = _T_90 ^ _T_91; // @[convert.scala 18:36]
  assign _T_93 = io_B[6:1]; // @[convert.scala 19:24]
  assign _T_94 = io_B[5:0]; // @[convert.scala 19:43]
  assign _T_95 = _T_93 ^ _T_94; // @[convert.scala 19:39]
  assign _T_96 = _T_95[5:2]; // @[LZD.scala 43:32]
  assign _T_97 = _T_96[3:2]; // @[LZD.scala 43:32]
  assign _T_98 = _T_97 != 2'h0; // @[LZD.scala 39:14]
  assign _T_99 = _T_97[1]; // @[LZD.scala 39:21]
  assign _T_100 = _T_97[0]; // @[LZD.scala 39:30]
  assign _T_101 = ~ _T_100; // @[LZD.scala 39:27]
  assign _T_102 = _T_99 | _T_101; // @[LZD.scala 39:25]
  assign _T_103 = {_T_98,_T_102}; // @[Cat.scala 29:58]
  assign _T_104 = _T_96[1:0]; // @[LZD.scala 44:32]
  assign _T_105 = _T_104 != 2'h0; // @[LZD.scala 39:14]
  assign _T_106 = _T_104[1]; // @[LZD.scala 39:21]
  assign _T_107 = _T_104[0]; // @[LZD.scala 39:30]
  assign _T_108 = ~ _T_107; // @[LZD.scala 39:27]
  assign _T_109 = _T_106 | _T_108; // @[LZD.scala 39:25]
  assign _T_110 = {_T_105,_T_109}; // @[Cat.scala 29:58]
  assign _T_111 = _T_103[1]; // @[Shift.scala 12:21]
  assign _T_112 = _T_110[1]; // @[Shift.scala 12:21]
  assign _T_113 = _T_111 | _T_112; // @[LZD.scala 49:16]
  assign _T_114 = ~ _T_112; // @[LZD.scala 49:27]
  assign _T_115 = _T_111 | _T_114; // @[LZD.scala 49:25]
  assign _T_116 = _T_103[0:0]; // @[LZD.scala 49:47]
  assign _T_117 = _T_110[0:0]; // @[LZD.scala 49:59]
  assign _T_118 = _T_111 ? _T_116 : _T_117; // @[LZD.scala 49:35]
  assign _T_120 = {_T_113,_T_115,_T_118}; // @[Cat.scala 29:58]
  assign _T_121 = _T_95[1:0]; // @[LZD.scala 44:32]
  assign _T_122 = _T_121 != 2'h0; // @[LZD.scala 39:14]
  assign _T_123 = _T_121[1]; // @[LZD.scala 39:21]
  assign _T_124 = _T_121[0]; // @[LZD.scala 39:30]
  assign _T_125 = ~ _T_124; // @[LZD.scala 39:27]
  assign _T_126 = _T_123 | _T_125; // @[LZD.scala 39:25]
  assign _T_127 = {_T_122,_T_126}; // @[Cat.scala 29:58]
  assign _T_128 = _T_120[2]; // @[Shift.scala 12:21]
  assign _T_130 = _T_120[1:0]; // @[LZD.scala 55:32]
  assign _T_131 = _T_128 ? _T_130 : _T_127; // @[LZD.scala 55:20]
  assign _T_132 = {_T_128,_T_131}; // @[Cat.scala 29:58]
  assign _T_133 = ~ _T_132; // @[convert.scala 21:22]
  assign _T_134 = io_B[4:0]; // @[convert.scala 22:36]
  assign _T_135 = _T_133 < 3'h5; // @[Shift.scala 16:24]
  assign _T_137 = _T_133[2]; // @[Shift.scala 12:21]
  assign _T_138 = _T_134[0:0]; // @[Shift.scala 64:52]
  assign _T_140 = {_T_138,4'h0}; // @[Cat.scala 29:58]
  assign _T_141 = _T_137 ? _T_140 : _T_134; // @[Shift.scala 64:27]
  assign _T_142 = _T_133[1:0]; // @[Shift.scala 66:70]
  assign _T_143 = _T_142[1]; // @[Shift.scala 12:21]
  assign _T_144 = _T_141[2:0]; // @[Shift.scala 64:52]
  assign _T_146 = {_T_144,2'h0}; // @[Cat.scala 29:58]
  assign _T_147 = _T_143 ? _T_146 : _T_141; // @[Shift.scala 64:27]
  assign _T_148 = _T_142[0:0]; // @[Shift.scala 66:70]
  assign _T_150 = _T_147[3:0]; // @[Shift.scala 64:52]
  assign _T_151 = {_T_150,1'h0}; // @[Cat.scala 29:58]
  assign _T_152 = _T_148 ? _T_151 : _T_147; // @[Shift.scala 64:27]
  assign _T_153 = _T_135 ? _T_152 : 5'h0; // @[Shift.scala 16:10]
  assign _T_154 = _T_153[4:4]; // @[convert.scala 23:34]
  assign decB_fraction = _T_153[3:0]; // @[convert.scala 24:34]
  assign _T_156 = _T_92 == 1'h0; // @[convert.scala 25:26]
  assign _T_158 = _T_92 ? _T_133 : _T_132; // @[convert.scala 25:42]
  assign _T_161 = ~ _T_154; // @[convert.scala 26:67]
  assign _T_162 = _T_90 ? _T_161 : _T_154; // @[convert.scala 26:51]
  assign _T_163 = {_T_156,_T_158,_T_162}; // @[Cat.scala 29:58]
  assign _T_165 = io_B[6:0]; // @[convert.scala 29:56]
  assign _T_166 = _T_165 != 7'h0; // @[convert.scala 29:60]
  assign _T_167 = ~ _T_166; // @[convert.scala 29:41]
  assign decB_isNaR = _T_90 & _T_167; // @[convert.scala 29:39]
  assign _T_170 = _T_90 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_170 & _T_167; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_163); // @[convert.scala 32:24]
  assign _T_178 = ~ _T_1; // @[PositMultiplier.scala 43:34]
  assign _T_180 = {_T_1,_T_178,decA_fraction}; // @[Cat.scala 29:58]
  assign sigA = $signed(_T_180); // @[PositMultiplier.scala 43:61]
  assign _T_181 = ~ _T_90; // @[PositMultiplier.scala 44:34]
  assign _T_183 = {_T_90,_T_181,decB_fraction}; // @[Cat.scala 29:58]
  assign sigB = $signed(_T_183); // @[PositMultiplier.scala 44:61]
  assign _T_184 = $signed(sigA) * $signed(sigB); // @[PositMultiplier.scala 45:25]
  assign sigP = $unsigned(_T_184); // @[PositMultiplier.scala 45:33]
  assign head2 = sigP[11:10]; // @[PositMultiplier.scala 46:28]
  assign _T_185 = head2[1]; // @[PositMultiplier.scala 47:31]
  assign _T_186 = ~ _T_185; // @[PositMultiplier.scala 47:25]
  assign _T_187 = head2[0]; // @[PositMultiplier.scala 47:42]
  assign addTwo = _T_186 & _T_187; // @[PositMultiplier.scala 47:35]
  assign _T_188 = sigP[11]; // @[PositMultiplier.scala 49:23]
  assign _T_189 = sigP[9]; // @[PositMultiplier.scala 49:49]
  assign addOne = _T_188 ^ _T_189; // @[PositMultiplier.scala 49:43]
  assign _T_190 = {addTwo,addOne}; // @[Cat.scala 29:58]
  assign expBias = {1'b0,$signed(_T_190)}; // @[PositMultiplier.scala 50:39]
  assign _T_191 = sigP[8:0]; // @[PositMultiplier.scala 53:81]
  assign _T_192 = sigP[7:0]; // @[PositMultiplier.scala 54:81]
  assign _T_193 = {_T_192, 1'h0}; // @[PositMultiplier.scala 54:104]
  assign frac = addOne ? _T_191 : _T_193; // @[PositMultiplier.scala 51:22]
  assign _T_194 = $signed(decA_scale) + $signed(decB_scale); // @[PositMultiplier.scala 56:30]
  assign _GEN_0 = {{3{expBias[2]}},expBias}; // @[PositMultiplier.scala 56:44]
  assign _T_196 = $signed(_T_194) + $signed(_GEN_0); // @[PositMultiplier.scala 56:44]
  assign mulScale = $signed(_T_196); // @[PositMultiplier.scala 56:44]
  assign underflow = $signed(mulScale) < $signed(-6'shd); // @[PositMultiplier.scala 57:28]
  assign overflow = $signed(mulScale) > $signed(6'shc); // @[PositMultiplier.scala 58:28]
  assign decM_sign = sigP[11:11]; // @[PositMultiplier.scala 62:29]
  assign _T_199 = underflow ? $signed(-6'shd) : $signed(mulScale); // @[Mux.scala 87:16]
  assign _T_200 = overflow ? $signed(6'shc) : $signed(_T_199); // @[Mux.scala 87:16]
  assign decM_fraction = frac[8:5]; // @[PositMultiplier.scala 70:29]
  assign decM_isNaR = decA_isNaR | decB_isNaR; // @[PositMultiplier.scala 71:31]
  assign decM_isZero = decA_isZero | decB_isZero; // @[PositMultiplier.scala 72:32]
  assign grsTmp = frac[4:0]; // @[PositMultiplier.scala 75:30]
  assign _T_204 = grsTmp[4:3]; // @[PositMultiplier.scala 78:32]
  assign _T_205 = grsTmp[2:0]; // @[PositMultiplier.scala 78:48]
  assign _T_206 = _T_205 != 3'h0; // @[PositMultiplier.scala 78:52]
  assign _GEN_1 = _T_200[4:0]; // @[PositMultiplier.scala 60:23 PositMultiplier.scala 63:17]
  assign decM_scale = $signed(_GEN_1); // @[PositMultiplier.scala 60:23 PositMultiplier.scala 63:17]
  assign _T_209 = decM_scale[0]; // @[convert.scala 46:61]
  assign _T_210 = ~ _T_209; // @[convert.scala 46:52]
  assign _T_212 = decM_sign ? _T_210 : _T_209; // @[convert.scala 46:42]
  assign _T_213 = decM_scale[4:1]; // @[convert.scala 48:34]
  assign _T_214 = _T_213[3:3]; // @[convert.scala 49:36]
  assign _T_216 = ~ _T_213; // @[convert.scala 50:36]
  assign _T_217 = $signed(_T_216); // @[convert.scala 50:36]
  assign _T_218 = _T_214 ? $signed(_T_217) : $signed(_T_213); // @[convert.scala 50:28]
  assign _T_219 = _T_214 ^ decM_sign; // @[convert.scala 51:31]
  assign _T_220 = ~ _T_219; // @[convert.scala 52:43]
  assign _T_224 = {_T_220,_T_219,_T_212,decM_fraction,_T_204,_T_206}; // @[Cat.scala 29:58]
  assign _T_225 = $unsigned(_T_218); // @[Shift.scala 39:17]
  assign _T_226 = _T_225 < 4'ha; // @[Shift.scala 39:24]
  assign _T_228 = _T_224[9:8]; // @[Shift.scala 90:30]
  assign _T_229 = _T_224[7:0]; // @[Shift.scala 90:48]
  assign _T_230 = _T_229 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_2 = {{1'd0}, _T_230}; // @[Shift.scala 90:39]
  assign _T_231 = _T_228 | _GEN_2; // @[Shift.scala 90:39]
  assign _T_232 = _T_225[3]; // @[Shift.scala 12:21]
  assign _T_233 = _T_224[9]; // @[Shift.scala 12:21]
  assign _T_235 = _T_233 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_236 = {_T_235,_T_231}; // @[Cat.scala 29:58]
  assign _T_237 = _T_232 ? _T_236 : _T_224; // @[Shift.scala 91:22]
  assign _T_238 = _T_225[2:0]; // @[Shift.scala 92:77]
  assign _T_239 = _T_237[9:4]; // @[Shift.scala 90:30]
  assign _T_240 = _T_237[3:0]; // @[Shift.scala 90:48]
  assign _T_241 = _T_240 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_3 = {{5'd0}, _T_241}; // @[Shift.scala 90:39]
  assign _T_242 = _T_239 | _GEN_3; // @[Shift.scala 90:39]
  assign _T_243 = _T_238[2]; // @[Shift.scala 12:21]
  assign _T_244 = _T_237[9]; // @[Shift.scala 12:21]
  assign _T_246 = _T_244 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_247 = {_T_246,_T_242}; // @[Cat.scala 29:58]
  assign _T_248 = _T_243 ? _T_247 : _T_237; // @[Shift.scala 91:22]
  assign _T_249 = _T_238[1:0]; // @[Shift.scala 92:77]
  assign _T_250 = _T_248[9:2]; // @[Shift.scala 90:30]
  assign _T_251 = _T_248[1:0]; // @[Shift.scala 90:48]
  assign _T_252 = _T_251 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_4 = {{7'd0}, _T_252}; // @[Shift.scala 90:39]
  assign _T_253 = _T_250 | _GEN_4; // @[Shift.scala 90:39]
  assign _T_254 = _T_249[1]; // @[Shift.scala 12:21]
  assign _T_255 = _T_248[9]; // @[Shift.scala 12:21]
  assign _T_257 = _T_255 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_258 = {_T_257,_T_253}; // @[Cat.scala 29:58]
  assign _T_259 = _T_254 ? _T_258 : _T_248; // @[Shift.scala 91:22]
  assign _T_260 = _T_249[0:0]; // @[Shift.scala 92:77]
  assign _T_261 = _T_259[9:1]; // @[Shift.scala 90:30]
  assign _T_262 = _T_259[0:0]; // @[Shift.scala 90:48]
  assign _GEN_5 = {{8'd0}, _T_262}; // @[Shift.scala 90:39]
  assign _T_264 = _T_261 | _GEN_5; // @[Shift.scala 90:39]
  assign _T_266 = _T_259[9]; // @[Shift.scala 12:21]
  assign _T_267 = {_T_266,_T_264}; // @[Cat.scala 29:58]
  assign _T_268 = _T_260 ? _T_267 : _T_259; // @[Shift.scala 91:22]
  assign _T_271 = _T_233 ? 10'h3ff : 10'h0; // @[Bitwise.scala 71:12]
  assign _T_272 = _T_226 ? _T_268 : _T_271; // @[Shift.scala 39:10]
  assign _T_273 = _T_272[3]; // @[convert.scala 55:31]
  assign _T_274 = _T_272[2]; // @[convert.scala 56:31]
  assign _T_275 = _T_272[1]; // @[convert.scala 57:31]
  assign _T_276 = _T_272[0]; // @[convert.scala 58:31]
  assign _T_277 = _T_272[9:3]; // @[convert.scala 59:69]
  assign _T_278 = _T_277 != 7'h0; // @[convert.scala 59:81]
  assign _T_279 = ~ _T_278; // @[convert.scala 59:50]
  assign _T_281 = _T_277 == 7'h7f; // @[convert.scala 60:81]
  assign _T_282 = _T_273 | _T_275; // @[convert.scala 61:44]
  assign _T_283 = _T_282 | _T_276; // @[convert.scala 61:52]
  assign _T_284 = _T_274 & _T_283; // @[convert.scala 61:36]
  assign _T_285 = ~ _T_281; // @[convert.scala 62:63]
  assign _T_286 = _T_285 & _T_284; // @[convert.scala 62:103]
  assign _T_287 = _T_279 | _T_286; // @[convert.scala 62:60]
  assign _GEN_6 = {{6'd0}, _T_287}; // @[convert.scala 63:56]
  assign _T_290 = _T_277 + _GEN_6; // @[convert.scala 63:56]
  assign _T_291 = {decM_sign,_T_290}; // @[Cat.scala 29:58]
  assign _T_293 = decM_isZero ? 8'h0 : _T_291; // @[Mux.scala 87:16]
  assign io_M = decM_isNaR ? 8'h80 : _T_293; // @[PositMultiplier.scala 86:8]
endmodule
